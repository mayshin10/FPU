
module FPU_normalize ( src, result, shifted );
  input [24:0] src;
  output [22:0] result;
  output [4:0] shifted;
  wire   n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n92, n93, n94, n95,
         n1, n2, n4, n5, n18, n28, n63, n90, n91, n97, n99, n101;

  AND3X1_RVT U113 ( .A1(shifted[4]), .A2(n69), .A3(src[0]), .Y(n68) );
  NOR4X0_RVT U114 ( .A1(n44), .A2(n36), .A3(n83), .A4(n81), .Y(shifted[2]) );
  OR4X1_RVT U118 ( .A1(src[18]), .A2(src[19]), .A3(src[20]), .A4(src[21]), .Y(
        n95) );
  OR4X1_RVT U119 ( .A1(src[22]), .A2(src[23]), .A3(src[24]), .A4(src[9]), .Y(
        n94) );
  OR4X1_RVT U120 ( .A1(src[10]), .A2(src[11]), .A3(src[12]), .A4(src[13]), .Y(
        n93) );
  OR4X1_RVT U121 ( .A1(src[14]), .A2(src[15]), .A3(src[16]), .A4(src[17]), .Y(
        n92) );
  AO22X1_RVT U2 ( .A1(shifted[0]), .A2(n31), .A3(n32), .A4(n91), .Y(result[22]) );
  AO22X1_RVT U3 ( .A1(n57), .A2(n90), .A3(shifted[0]), .A4(n60), .Y(result[16]) );
  AO22X1_RVT U4 ( .A1(n54), .A2(n91), .A3(shifted[0]), .A4(n57), .Y(result[17]) );
  AO22X1_RVT U5 ( .A1(n51), .A2(n91), .A3(shifted[0]), .A4(n54), .Y(result[18]) );
  AO22X1_RVT U6 ( .A1(n46), .A2(n91), .A3(shifted[0]), .A4(n51), .Y(result[19]) );
  AO22X1_RVT U7 ( .A1(n31), .A2(n91), .A3(shifted[0]), .A4(n38), .Y(result[21]) );
  AOI221X1_RVT U8 ( .A1(n33), .A2(n41), .A3(n35), .A4(n44), .A5(n79), .Y(n1)
         );
  AND2X1_RVT U9 ( .A1(n69), .A2(n101), .Y(n2) );
  NOR4X0_RVT U10 ( .A1(n92), .A2(n93), .A3(n94), .A4(n95), .Y(shifted[4]) );
  AND2X1_RVT U11 ( .A1(shifted[1]), .A2(n91), .Y(n14) );
  AND2X1_RVT U12 ( .A1(n43), .A2(n2), .Y(n30) );
  AND2X1_RVT U13 ( .A1(n2), .A2(n35), .Y(n26) );
  INVX1_RVT U14 ( .A(n1), .Y(n91) );
  INVX1_RVT U15 ( .A(n4), .Y(n63) );
  INVX1_RVT U16 ( .A(n4), .Y(n28) );
  INVX1_RVT U17 ( .A(n12), .Y(shifted[1]) );
  AND2X1_RVT U18 ( .A1(shifted[1]), .A2(n99), .Y(n35) );
  AND2X1_RVT U19 ( .A1(n12), .A2(n99), .Y(n43) );
  INVX1_RVT U20 ( .A(shifted[0]), .Y(n90) );
  AND2X1_RVT U21 ( .A1(n91), .A2(n12), .Y(n6) );
  AND2X1_RVT U22 ( .A1(n2), .A2(n99), .Y(n23) );
  AND2X1_RVT U23 ( .A1(shifted[0]), .A2(shifted[1]), .Y(n16) );
  AND2X1_RVT U24 ( .A1(shifted[0]), .A2(n12), .Y(n8) );
  NAND2X0_RVT U25 ( .A1(shifted[3]), .A2(n101), .Y(n4) );
  AND2X1_RVT U26 ( .A1(shifted[1]), .A2(shifted[2]), .Y(n33) );
  OR2X1_RVT U27 ( .A1(n37), .A2(n79), .Y(n12) );
  INVX1_RVT U28 ( .A(shifted[2]), .Y(n99) );
  INVX1_RVT U29 ( .A(n69), .Y(shifted[3]) );
  INVX1_RVT U30 ( .A(n97), .Y(shifted[0]) );
  INVX1_RVT U31 ( .A(n1), .Y(n97) );
  AND2X1_RVT U32 ( .A1(shifted[2]), .A2(n12), .Y(n40) );
  AO22X1_RVT U33 ( .A1(n38), .A2(n91), .A3(shifted[0]), .A4(n46), .Y(
        result[20]) );
  AO22X1_RVT U34 ( .A1(n60), .A2(n90), .A3(shifted[0]), .A4(n65), .Y(
        result[15]) );
  AO22X1_RVT U35 ( .A1(n70), .A2(n91), .A3(shifted[0]), .A4(n73), .Y(
        result[13]) );
  AO22X1_RVT U36 ( .A1(n65), .A2(n91), .A3(shifted[0]), .A4(n70), .Y(
        result[14]) );
  AO22X1_RVT U37 ( .A1(n73), .A2(n90), .A3(shifted[0]), .A4(n76), .Y(
        result[12]) );
  AO22X1_RVT U38 ( .A1(n11), .A2(n12), .A3(shifted[1]), .A4(n13), .Y(result[8]) );
  AND2X1_RVT U39 ( .A1(n2), .A2(shifted[2]), .Y(n22) );
  AO221X1_RVT U40 ( .A1(n33), .A2(n34), .A3(n35), .A4(n36), .A5(n37), .Y(n32)
         );
  INVX1_RVT U41 ( .A(shifted[4]), .Y(n101) );
  AO21X1_RVT U42 ( .A1(shifted[2]), .A2(n45), .A3(n81), .Y(n79) );
  AO21X1_RVT U43 ( .A1(shifted[2]), .A2(n49), .A3(n83), .Y(n37) );
  NAND2X0_RVT U44 ( .A1(n5), .A2(n18), .Y(n69) );
  NOR4X1_RVT U45 ( .A1(n88), .A2(n89), .A3(n87), .A4(n86), .Y(n5) );
  NOR4X1_RVT U46 ( .A1(n64), .A2(n80), .A3(n84), .A4(n82), .Y(n18) );
  AO221X1_RVT U47 ( .A1(n33), .A2(n61), .A3(n40), .A4(n55), .A5(n62), .Y(n57)
         );
  AO22X1_RVT U48 ( .A1(n43), .A2(n34), .A3(n35), .A4(n47), .Y(n62) );
  AO221X1_RVT U49 ( .A1(n33), .A2(n66), .A3(n40), .A4(n58), .A5(n67), .Y(n60)
         );
  AO22X1_RVT U50 ( .A1(n43), .A2(n39), .A3(n35), .A4(n52), .Y(n67) );
  AO221X1_RVT U51 ( .A1(n33), .A2(n58), .A3(n40), .A4(n52), .A5(n59), .Y(n54)
         );
  AO22X1_RVT U52 ( .A1(n43), .A2(n41), .A3(n35), .A4(n39), .Y(n59) );
  AO221X1_RVT U53 ( .A1(n33), .A2(n47), .A3(n40), .A4(n34), .A5(n48), .Y(n38)
         );
  AO22X1_RVT U54 ( .A1(n43), .A2(n36), .A3(n35), .A4(n49), .Y(n48) );
  AO221X1_RVT U55 ( .A1(n33), .A2(n52), .A3(n40), .A4(n39), .A5(n53), .Y(n46)
         );
  AO22X1_RVT U56 ( .A1(n43), .A2(n45), .A3(n35), .A4(n41), .Y(n53) );
  AO221X1_RVT U57 ( .A1(n33), .A2(n55), .A3(n40), .A4(n47), .A5(n56), .Y(n51)
         );
  AO22X1_RVT U58 ( .A1(n43), .A2(n49), .A3(n35), .A4(n34), .Y(n56) );
  AO221X1_RVT U59 ( .A1(n33), .A2(n39), .A3(n40), .A4(n41), .A5(n42), .Y(n31)
         );
  AO22X1_RVT U60 ( .A1(n43), .A2(n44), .A3(n35), .A4(n45), .Y(n42) );
  AO221X1_RVT U61 ( .A1(n33), .A2(n71), .A3(n40), .A4(n61), .A5(n72), .Y(n65)
         );
  AO22X1_RVT U62 ( .A1(n43), .A2(n47), .A3(n35), .A4(n55), .Y(n72) );
  AO22X1_RVT U63 ( .A1(n24), .A2(n91), .A3(shifted[0]), .A4(n25), .Y(result[4]) );
  AO22X1_RVT U64 ( .A1(n29), .A2(n90), .A3(n50), .A4(n30), .Y(result[1]) );
  AO22X1_RVT U65 ( .A1(n90), .A2(n20), .A3(shifted[0]), .A4(n15), .Y(n13) );
  AO22X1_RVT U66 ( .A1(n90), .A2(n9), .A3(shifted[0]), .A4(n19), .Y(n11) );
  AO22X1_RVT U67 ( .A1(n27), .A2(n91), .A3(shifted[0]), .A4(n29), .Y(result[2]) );
  AO22X1_RVT U68 ( .A1(n25), .A2(n91), .A3(shifted[0]), .A4(n27), .Y(result[3]) );
  AO22X1_RVT U69 ( .A1(n91), .A2(n19), .A3(shifted[0]), .A4(n20), .Y(n10) );
  AO222X1_RVT U70 ( .A1(n6), .A2(n77), .A3(n8), .A4(n7), .A5(shifted[1]), .A6(
        n11), .Y(result[10]) );
  AO222X1_RVT U71 ( .A1(n14), .A2(n17), .A3(n16), .A4(n21), .A5(n13), .A6(n12), 
        .Y(result[6]) );
  AO222X1_RVT U72 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .A5(shifted[1]), .A6(
        n10), .Y(result[9]) );
  AO222X1_RVT U73 ( .A1(n6), .A2(n15), .A3(n14), .A4(n21), .A5(shifted[0]), 
        .A6(n24), .Y(result[5]) );
  AO222X1_RVT U74 ( .A1(n14), .A2(n15), .A3(n16), .A4(n17), .A5(n10), .A6(n12), 
        .Y(result[7]) );
  AO222X1_RVT U75 ( .A1(n8), .A2(n77), .A3(n16), .A4(n9), .A5(n76), .A6(n91), 
        .Y(result[11]) );
  AND2X1_RVT U76 ( .A1(n30), .A2(n78), .Y(result[0]) );
  AO222X1_RVT U77 ( .A1(n43), .A2(n58), .A3(n40), .A4(n74), .A5(shifted[1]), 
        .A6(n7), .Y(n76) );
  AO222X1_RVT U78 ( .A1(n43), .A2(n55), .A3(n40), .A4(n71), .A5(shifted[1]), 
        .A6(n77), .Y(n73) );
  AO221X1_RVT U79 ( .A1(n33), .A2(n74), .A3(n40), .A4(n66), .A5(n75), .Y(n70)
         );
  AO22X1_RVT U80 ( .A1(n43), .A2(n52), .A3(n35), .A4(n58), .Y(n75) );
  AO221X1_RVT U81 ( .A1(n85), .A2(src[0]), .A3(src[16]), .A4(n28), .A5(n86), 
        .Y(n81) );
  AND2X1_RVT U82 ( .A1(shifted[3]), .A2(shifted[4]), .Y(n85) );
  AO21X1_RVT U83 ( .A1(src[10]), .A2(n63), .A3(n80), .Y(n41) );
  AO21X1_RVT U84 ( .A1(src[13]), .A2(n63), .A3(n88), .Y(n36) );
  AO21X1_RVT U85 ( .A1(src[14]), .A2(n63), .A3(n89), .Y(n44) );
  AO21X1_RVT U86 ( .A1(src[12]), .A2(n63), .A3(n82), .Y(n45) );
  AO21X1_RVT U87 ( .A1(src[15]), .A2(n63), .A3(n87), .Y(n83) );
  AO21X1_RVT U88 ( .A1(src[8]), .A2(shifted[4]), .A3(src[24]), .Y(n86) );
  AO21X1_RVT U89 ( .A1(src[4]), .A2(shifted[4]), .A3(src[20]), .Y(n82) );
  AO21X1_RVT U90 ( .A1(src[7]), .A2(shifted[4]), .A3(src[23]), .Y(n87) );
  AO21X1_RVT U91 ( .A1(src[3]), .A2(shifted[4]), .A3(src[19]), .Y(n84) );
  AO21X1_RVT U92 ( .A1(src[6]), .A2(shifted[4]), .A3(src[22]), .Y(n89) );
  AO21X1_RVT U93 ( .A1(src[2]), .A2(shifted[4]), .A3(src[18]), .Y(n80) );
  AO21X1_RVT U94 ( .A1(src[5]), .A2(shifted[4]), .A3(src[21]), .Y(n88) );
  AO21X1_RVT U95 ( .A1(src[1]), .A2(shifted[4]), .A3(src[17]), .Y(n64) );
  AO21X1_RVT U96 ( .A1(src[11]), .A2(n63), .A3(n84), .Y(n49) );
  AO22X1_RVT U97 ( .A1(n2), .A2(src[13]), .A3(n28), .A4(src[5]), .Y(n55) );
  AO22X1_RVT U98 ( .A1(n2), .A2(src[12]), .A3(n28), .A4(src[4]), .Y(n58) );
  AO22X1_RVT U99 ( .A1(n2), .A2(src[15]), .A3(n63), .A4(src[7]), .Y(n47) );
  AO22X1_RVT U100 ( .A1(n2), .A2(src[14]), .A3(n63), .A4(src[6]), .Y(n52) );
  AO22X1_RVT U101 ( .A1(n2), .A2(src[10]), .A3(n28), .A4(src[2]), .Y(n66) );
  AO22X1_RVT U102 ( .A1(n2), .A2(src[11]), .A3(n28), .A4(src[3]), .Y(n61) );
  AO21X1_RVT U103 ( .A1(src[9]), .A2(n63), .A3(n64), .Y(n34) );
  AO221X1_RVT U104 ( .A1(n28), .A2(src[8]), .A3(n2), .A4(src[16]), .A5(n68), 
        .Y(n39) );
  AO22X1_RVT U105 ( .A1(src[9]), .A2(n2), .A3(n28), .A4(src[1]), .Y(n71) );
  AO22X1_RVT U106 ( .A1(src[1]), .A2(n91), .A3(shifted[0]), .A4(src[0]), .Y(
        n78) );
  AO22X1_RVT U107 ( .A1(n2), .A2(src[8]), .A3(n28), .A4(src[0]), .Y(n74) );
  AO22X1_RVT U108 ( .A1(n61), .A2(n99), .A3(n22), .A4(src[7]), .Y(n77) );
  AO22X1_RVT U109 ( .A1(n99), .A2(n66), .A3(n22), .A4(src[6]), .Y(n7) );
  AO22X1_RVT U110 ( .A1(n71), .A2(n99), .A3(n22), .A4(src[5]), .Y(n9) );
  AO22X1_RVT U111 ( .A1(n22), .A2(src[2]), .A3(n23), .A4(src[6]), .Y(n15) );
  AO22X1_RVT U112 ( .A1(n22), .A2(src[1]), .A3(n23), .A4(src[5]), .Y(n17) );
  AO22X1_RVT U115 ( .A1(n22), .A2(src[0]), .A3(n23), .A4(src[4]), .Y(n21) );
  AO22X1_RVT U116 ( .A1(n74), .A2(n99), .A3(n22), .A4(src[4]), .Y(n19) );
  AO22X1_RVT U117 ( .A1(n17), .A2(n12), .A3(n26), .A4(src[3]), .Y(n24) );
  AO22X1_RVT U122 ( .A1(n22), .A2(src[3]), .A3(n23), .A4(src[7]), .Y(n20) );
  AO22X1_RVT U123 ( .A1(n30), .A2(src[2]), .A3(n26), .A4(src[0]), .Y(n29) );
  AO22X1_RVT U124 ( .A1(n30), .A2(src[3]), .A3(n26), .A4(src[1]), .Y(n27) );
  AO22X1_RVT U125 ( .A1(n21), .A2(n12), .A3(n26), .A4(src[2]), .Y(n25) );
  AND2X1_RVT U126 ( .A1(shifted[0]), .A2(src[1]), .Y(n50) );
endmodule


module FPU_CAL_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HADDX1_RVT U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1_RVT U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1_RVT U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1_RVT U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1_RVT U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1_RVT U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX1_RVT U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1_RVT U2 ( .A1(carry[7]), .A2(A[7]), .Y(SUM[7]) );
endmodule


module FPU_CAL_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HADDX1_RVT U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1_RVT U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1_RVT U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1_RVT U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1_RVT U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1_RVT U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX1_RVT U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1_RVT U2 ( .A1(carry[7]), .A2(A[7]), .Y(SUM[7]) );
endmodule


module FPU_CAL_DW01_inc_2 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HADDX1_RVT U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1_RVT U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1_RVT U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1_RVT U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1_RVT U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1_RVT U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX1_RVT U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1_RVT U2 ( .A1(carry[7]), .A2(A[7]), .Y(SUM[7]) );
endmodule


module FPU_CAL_DW01_inc_3 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1_RVT U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1_RVT U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1_RVT U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1_RVT U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1_RVT U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1_RVT U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1_RVT U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX1_RVT U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1_RVT U2 ( .A1(carry[8]), .A2(A[8]), .Y(SUM[8]) );
endmodule


module FPU_CAL_DW01_add_0 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .S(SUM[7])
         );
  AND2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
  XOR2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
endmodule


module FPU_CAL_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] DIFF;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [25:0] carry;

  FADDX1_RVT U2_13 ( .A(A[13]), .B(n6), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FADDX1_RVT U2_11 ( .A(A[11]), .B(n4), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FADDX1_RVT U2_12 ( .A(A[12]), .B(n5), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FADDX1_RVT U2_15 ( .A(A[15]), .B(n7), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FADDX1_RVT U2_16 ( .A(A[16]), .B(n15), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FADDX1_RVT U2_18 ( .A(A[18]), .B(n17), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FADDX1_RVT U2_19 ( .A(A[19]), .B(n18), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FADDX1_RVT U2_1 ( .A(A[1]), .B(n23), .CI(carry[1]), .CO(carry[2]), .S(
        DIFF[1]) );
  FADDX1_RVT U2_2 ( .A(A[2]), .B(n24), .CI(carry[2]), .CO(carry[3]), .S(
        DIFF[2]) );
  FADDX1_RVT U2_4 ( .A(A[4]), .B(n8), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FADDX1_RVT U2_9 ( .A(A[9]), .B(n14), .CI(carry[9]), .CO(carry[10]), .S(
        DIFF[9]) );
  FADDX1_RVT U2_3 ( .A(A[3]), .B(n25), .CI(carry[3]), .CO(carry[4]), .S(
        DIFF[3]) );
  FADDX1_RVT U2_7 ( .A(A[7]), .B(n11), .CI(carry[7]), .CO(carry[8]), .S(
        DIFF[7]) );
  FADDX1_RVT U2_6 ( .A(A[6]), .B(n10), .CI(carry[6]), .CO(carry[7]), .S(
        DIFF[6]) );
  FADDX1_RVT U2_5 ( .A(A[5]), .B(n9), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FADDX1_RVT U2_17 ( .A(A[17]), .B(n16), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FADDX1_RVT U2_21 ( .A(A[21]), .B(n21), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FADDX1_RVT U2_20 ( .A(A[20]), .B(n20), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FADDX1_RVT U2_22 ( .A(A[22]), .B(n19), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FADDX1_RVT U2_14 ( .A(A[14]), .B(n12), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FADDX1_RVT U2_10 ( .A(A[10]), .B(n3), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1_RVT U2_8 ( .A(A[8]), .B(n13), .CI(carry[8]), .CO(carry[9]), .S(
        DIFF[8]) );
  FADDX1_RVT U2_23 ( .A(A[23]), .B(n22), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  INVX1_RVT U1 ( .A(B[13]), .Y(n6) );
  XNOR2X1_RVT U2 ( .A1(A[0]), .A2(n2), .Y(DIFF[0]) );
  INVX1_RVT U3 ( .A(B[9]), .Y(n14) );
  INVX1_RVT U4 ( .A(B[17]), .Y(n16) );
  INVX1_RVT U5 ( .A(B[5]), .Y(n9) );
  INVX1_RVT U6 ( .A(B[6]), .Y(n10) );
  INVX1_RVT U7 ( .A(B[10]), .Y(n3) );
  INVX1_RVT U8 ( .A(B[12]), .Y(n5) );
  INVX1_RVT U9 ( .A(B[3]), .Y(n25) );
  INVX1_RVT U10 ( .A(B[7]), .Y(n11) );
  INVX0_RVT U11 ( .A(B[0]), .Y(n2) );
  INVX1_RVT U12 ( .A(B[8]), .Y(n13) );
  INVX0_RVT U13 ( .A(B[2]), .Y(n24) );
  INVX0_RVT U14 ( .A(B[4]), .Y(n8) );
  INVX1_RVT U15 ( .A(B[23]), .Y(n22) );
  INVX0_RVT U16 ( .A(B[11]), .Y(n4) );
  INVX0_RVT U17 ( .A(B[14]), .Y(n12) );
  INVX1_RVT U18 ( .A(B[18]), .Y(n17) );
  INVX1_RVT U19 ( .A(B[19]), .Y(n18) );
  INVX1_RVT U20 ( .A(B[15]), .Y(n7) );
  INVX1_RVT U21 ( .A(B[22]), .Y(n19) );
  INVX1_RVT U22 ( .A(B[20]), .Y(n20) );
  INVX1_RVT U23 ( .A(B[21]), .Y(n21) );
  INVX1_RVT U24 ( .A(B[16]), .Y(n15) );
  OR2X1_RVT U25 ( .A1(n2), .A2(A[0]), .Y(carry[1]) );
  INVX0_RVT U26 ( .A(B[1]), .Y(n23) );
  INVX1_RVT U27 ( .A(carry[24]), .Y(DIFF[24]) );
endmodule


module FPU_CAL_DW01_sub_3 ( A, B, CI, DIFF, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;
  wire   [25:0] carry;

  FADDX1_RVT U2_14 ( .A(A[14]), .B(n15), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FADDX1_RVT U2_15 ( .A(A[15]), .B(n10), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FADDX1_RVT U2_10 ( .A(A[10]), .B(n6), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1_RVT U2_11 ( .A(A[11]), .B(n7), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FADDX1_RVT U2_12 ( .A(A[12]), .B(n8), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FADDX1_RVT U2_7 ( .A(A[7]), .B(n14), .CI(carry[7]), .CO(carry[8]), .S(
        DIFF[7]) );
  FADDX1_RVT U2_8 ( .A(A[8]), .B(n16), .CI(carry[8]), .CO(carry[9]), .S(
        DIFF[8]) );
  FADDX1_RVT U2_3 ( .A(A[3]), .B(n28), .CI(carry[3]), .CO(carry[4]), .S(
        DIFF[3]) );
  FADDX1_RVT U2_1 ( .A(A[1]), .B(n26), .CI(carry[1]), .CO(carry[2]), .S(
        DIFF[1]) );
  FADDX1_RVT U2_5 ( .A(A[5]), .B(n12), .CI(carry[5]), .CO(carry[6]), .S(
        DIFF[5]) );
  FADDX1_RVT U2_6 ( .A(A[6]), .B(n13), .CI(carry[6]), .CO(carry[7]), .S(
        DIFF[6]) );
  FADDX1_RVT U2_2 ( .A(A[2]), .B(n27), .CI(carry[2]), .CO(carry[3]), .S(
        DIFF[2]) );
  FADDX1_RVT U2_21 ( .A(A[21]), .B(n24), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FADDX1_RVT U2_9 ( .A(A[9]), .B(n17), .CI(carry[9]), .CO(carry[10]), .S(
        DIFF[9]) );
  FADDX1_RVT U2_19 ( .A(A[19]), .B(n21), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FADDX1_RVT U2_18 ( .A(A[18]), .B(n20), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FADDX1_RVT U2_20 ( .A(A[20]), .B(n23), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FADDX1_RVT U2_22 ( .A(A[22]), .B(n22), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FADDX1_RVT U2_17 ( .A(A[17]), .B(n19), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FADDX1_RVT U2_16 ( .A(A[16]), .B(n18), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FADDX1_RVT U2_23 ( .A(A[23]), .B(n25), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  FADDX1_RVT U2_13 ( .A(A[13]), .B(n9), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  XNOR2X1_RVT U1 ( .A1(A[0]), .A2(n5), .Y(DIFF[0]) );
  NAND2X0_RVT U2 ( .A1(A[4]), .A2(carry[4]), .Y(n2) );
  NAND2X0_RVT U3 ( .A1(n11), .A2(carry[4]), .Y(n1) );
  XOR3X1_RVT U4 ( .A1(carry[4]), .A2(A[4]), .A3(n11), .Y(DIFF[4]) );
  NAND2X0_RVT U5 ( .A1(A[4]), .A2(n11), .Y(n3) );
  NAND3X0_RVT U6 ( .A1(n3), .A2(n2), .A3(n1), .Y(carry[5]) );
  INVX0_RVT U7 ( .A(B[23]), .Y(n25) );
  INVX0_RVT U8 ( .A(B[8]), .Y(n16) );
  INVX0_RVT U9 ( .A(B[5]), .Y(n12) );
  INVX0_RVT U10 ( .A(B[6]), .Y(n13) );
  INVX0_RVT U11 ( .A(B[7]), .Y(n14) );
  INVX0_RVT U12 ( .A(B[11]), .Y(n7) );
  INVX0_RVT U13 ( .A(B[15]), .Y(n10) );
  INVX1_RVT U14 ( .A(B[12]), .Y(n8) );
  INVX1_RVT U15 ( .A(B[16]), .Y(n18) );
  INVX1_RVT U16 ( .A(B[17]), .Y(n19) );
  INVX1_RVT U17 ( .A(B[22]), .Y(n22) );
  INVX1_RVT U18 ( .A(B[20]), .Y(n23) );
  INVX1_RVT U19 ( .A(B[18]), .Y(n20) );
  INVX1_RVT U20 ( .A(B[19]), .Y(n21) );
  INVX0_RVT U21 ( .A(B[13]), .Y(n9) );
  INVX0_RVT U22 ( .A(B[10]), .Y(n6) );
  INVX0_RVT U23 ( .A(B[9]), .Y(n17) );
  INVX1_RVT U24 ( .A(B[21]), .Y(n24) );
  INVX0_RVT U25 ( .A(B[14]), .Y(n15) );
  INVX0_RVT U26 ( .A(B[1]), .Y(n26) );
  OR2X1_RVT U27 ( .A1(n5), .A2(A[0]), .Y(carry[1]) );
  INVX0_RVT U28 ( .A(B[2]), .Y(n27) );
  INVX0_RVT U29 ( .A(B[3]), .Y(n28) );
  INVX1_RVT U30 ( .A(B[4]), .Y(n11) );
  INVX1_RVT U31 ( .A(B[0]), .Y(n5) );
  INVX1_RVT U32 ( .A(carry[24]), .Y(DIFF[24]) );
endmodule


module FPU_CAL_DW01_add_1 ( A, B, CI, SUM, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  input CI;
  output CO;

  wire   [24:1] carry;

  FADDX1_RVT U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1_RVT U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  FADDX1_RVT U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1_RVT U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1_RVT U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1_RVT U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  FADDX1_RVT U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1_RVT U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1_RVT U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1_RVT U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1_RVT U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1_RVT U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1_RVT U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1_RVT U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(SUM[24]), .S(
        SUM[23]) );
  AND2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
  XOR2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
endmodule


module FPU_CAL_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [23:0] A;
  input [7:0] SH;
  output [23:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117;

  INVX1_RVT U3 ( .A(SH[7]), .Y(n37) );
  INVX1_RVT U4 ( .A(n10), .Y(n77) );
  INVX1_RVT U5 ( .A(n25), .Y(n11) );
  NAND3X0_RVT U6 ( .A1(n12), .A2(n13), .A3(n5), .Y(n72) );
  NAND2X0_RVT U7 ( .A1(A[17]), .A2(n27), .Y(n8) );
  AO221X1_RVT U8 ( .A1(A[9]), .A2(n26), .A3(A[8]), .A4(n35), .A5(n113), .Y(n48) );
  AO22X1_RVT U9 ( .A1(A[11]), .A2(n34), .A3(A[10]), .A4(n31), .Y(n113) );
  NAND3X0_RVT U10 ( .A1(n14), .A2(n15), .A3(n16), .Y(B[12]) );
  INVX1_RVT U11 ( .A(n23), .Y(n36) );
  NAND2X0_RVT U12 ( .A1(SH[0]), .A2(SH[1]), .Y(n1) );
  AND2X1_RVT U13 ( .A1(n81), .A2(n98), .Y(n2) );
  OAI22X1_RVT U14 ( .A1(n20), .A2(n1), .A3(n21), .A4(n22), .Y(n3) );
  AO221X1_RVT U15 ( .A1(A[3]), .A2(n27), .A3(A[2]), .A4(n36), .A5(n3), .Y(n4)
         );
  AOI21X1_RVT U16 ( .A1(n36), .A2(A[20]), .A3(n33), .Y(n5) );
  AO22X1_RVT U17 ( .A1(n34), .A2(A[22]), .A3(n32), .A4(A[21]), .Y(n6) );
  AOI22X1_RVT U18 ( .A1(n33), .A2(A[19]), .A3(A[18]), .A4(n29), .Y(n7) );
  MUX21X1_RVT U19 ( .A1(n23), .A2(n11), .S0(n40), .Y(n10) );
  NAND2X0_RVT U20 ( .A1(A[16]), .A2(n35), .Y(n9) );
  NAND3X0_RVT U21 ( .A1(n8), .A2(n9), .A3(n7), .Y(n71) );
  NAND2X0_RVT U22 ( .A1(A[21]), .A2(SH[0]), .Y(n12) );
  NAND2X0_RVT U23 ( .A1(A[22]), .A2(SH[1]), .Y(n13) );
  NAND2X0_RVT U24 ( .A1(n43), .A2(n50), .Y(n14) );
  NAND2X0_RVT U25 ( .A1(n56), .A2(n72), .Y(n15) );
  NAND2X0_RVT U26 ( .A1(n2), .A2(n71), .Y(n16) );
  INVX1_RVT U27 ( .A(n88), .Y(n38) );
  INVX1_RVT U28 ( .A(n108), .Y(n39) );
  INVX1_RVT U29 ( .A(SH[0]), .Y(n42) );
  NAND2X0_RVT U30 ( .A1(n75), .A2(n4), .Y(n17) );
  NAND2X0_RVT U31 ( .A1(n73), .A2(n85), .Y(n18) );
  NAND3X0_RVT U32 ( .A1(n17), .A2(n18), .A3(n19), .Y(n84) );
  NAND2X0_RVT U33 ( .A1(n38), .A2(n86), .Y(n19) );
  INVX1_RVT U34 ( .A(A[4]), .Y(n21) );
  INVX1_RVT U35 ( .A(A[5]), .Y(n20) );
  NAND2X0_RVT U36 ( .A1(n42), .A2(SH[1]), .Y(n22) );
  INVX1_RVT U37 ( .A(n24), .Y(n26) );
  INVX1_RVT U38 ( .A(n22), .Y(n31) );
  INVX0_RVT U39 ( .A(n1), .Y(n34) );
  INVX1_RVT U40 ( .A(n1), .Y(n33) );
  NAND2X0_RVT U41 ( .A1(n42), .A2(n41), .Y(n23) );
  INVX1_RVT U42 ( .A(n24), .Y(n27) );
  INVX1_RVT U43 ( .A(n24), .Y(n28) );
  INVX1_RVT U44 ( .A(n22), .Y(n30) );
  INVX1_RVT U45 ( .A(n22), .Y(n32) );
  NAND2X0_RVT U46 ( .A1(SH[0]), .A2(n41), .Y(n24) );
  INVX1_RVT U47 ( .A(SH[1]), .Y(n41) );
  INVX1_RVT U48 ( .A(SH[2]), .Y(n40) );
  AO221X1_RVT U49 ( .A1(A[20]), .A2(n28), .A3(n35), .A4(A[19]), .A5(n6), .Y(
        n25) );
  AO221X1_RVT U50 ( .A1(A[16]), .A2(n28), .A3(A[15]), .A4(n35), .A5(n103), .Y(
        n57) );
  AND2X1_RVT U51 ( .A1(n84), .A2(n37), .Y(B[2]) );
  AO221X1_RVT U52 ( .A1(n43), .A2(n51), .A3(n2), .A4(n52), .A5(n53), .Y(B[7])
         );
  INVX1_RVT U53 ( .A(n23), .Y(n35) );
  AND2X1_RVT U54 ( .A1(n75), .A2(n37), .Y(n43) );
  AND2X1_RVT U55 ( .A1(n42), .A2(SH[1]), .Y(n29) );
  AO222X1_RVT U56 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .A5(n2), .A6(n47), 
        .Y(B[9]) );
  AO222X1_RVT U57 ( .A1(n43), .A2(n48), .A3(n45), .A4(n49), .A5(n2), .A6(n50), 
        .Y(B[8]) );
  AO222X1_RVT U58 ( .A1(n54), .A2(n25), .A3(n55), .A4(n35), .A5(n56), .A6(n57), 
        .Y(n53) );
  AO221X1_RVT U59 ( .A1(n43), .A2(n58), .A3(n2), .A4(n59), .A5(n60), .Y(B[6])
         );
  AO222X1_RVT U60 ( .A1(n56), .A2(n61), .A3(n54), .A4(n62), .A5(n63), .A6(n64), 
        .Y(n60) );
  AO221X1_RVT U61 ( .A1(n43), .A2(n65), .A3(n2), .A4(n44), .A5(n66), .Y(B[5])
         );
  AO222X1_RVT U62 ( .A1(n54), .A2(n67), .A3(n55), .A4(n68), .A5(n56), .A6(n47), 
        .Y(n66) );
  AO221X1_RVT U63 ( .A1(n43), .A2(n69), .A3(n2), .A4(n48), .A5(n70), .Y(B[4])
         );
  AO222X1_RVT U64 ( .A1(n54), .A2(n71), .A3(n55), .A4(n72), .A5(n56), .A6(n50), 
        .Y(n70) );
  AND2X1_RVT U65 ( .A1(n64), .A2(n40), .Y(n55) );
  AND2X1_RVT U66 ( .A1(n73), .A2(n37), .Y(n64) );
  AND2X1_RVT U67 ( .A1(n45), .A2(SH[2]), .Y(n54) );
  AND2X1_RVT U68 ( .A1(n74), .A2(n37), .Y(B[3]) );
  AO222X1_RVT U69 ( .A1(n75), .A2(n76), .A3(n73), .A4(n77), .A5(n38), .A6(n78), 
        .Y(n74) );
  AO222X1_RVT U70 ( .A1(n79), .A2(n57), .A3(n80), .A4(n52), .A5(n81), .A6(n51), 
        .Y(n78) );
  AO221X1_RVT U71 ( .A1(A[8]), .A2(n26), .A3(A[7]), .A4(n35), .A5(n82), .Y(n51) );
  AO22X1_RVT U72 ( .A1(A[10]), .A2(n34), .A3(A[9]), .A4(n30), .Y(n82) );
  AO221X1_RVT U73 ( .A1(A[4]), .A2(n28), .A3(A[3]), .A4(n36), .A5(n83), .Y(n76) );
  AO22X1_RVT U74 ( .A1(A[6]), .A2(n34), .A3(A[5]), .A4(n30), .Y(n83) );
  AO222X1_RVT U75 ( .A1(n79), .A2(n61), .A3(n80), .A4(n59), .A5(n81), .A6(n58), 
        .Y(n86) );
  AO221X1_RVT U76 ( .A1(A[7]), .A2(n28), .A3(A[6]), .A4(n36), .A5(n87), .Y(n58) );
  AO22X1_RVT U77 ( .A1(A[9]), .A2(n33), .A3(A[8]), .A4(n32), .Y(n87) );
  AND2X1_RVT U78 ( .A1(n39), .A2(n88), .Y(n73) );
  AND2X1_RVT U79 ( .A1(n43), .A2(n36), .Y(B[23]) );
  AND2X1_RVT U80 ( .A1(n89), .A2(n63), .Y(B[22]) );
  AND2X1_RVT U81 ( .A1(n43), .A2(n68), .Y(B[21]) );
  AND2X1_RVT U82 ( .A1(n43), .A2(n72), .Y(B[20]) );
  OA21X1_RVT U83 ( .A1(n90), .A2(n91), .A3(n37), .Y(B[1]) );
  MUX21X1_RVT U84 ( .A1(n92), .A2(n93), .S0(n38), .Y(n91) );
  AO222X1_RVT U85 ( .A1(n79), .A2(n47), .A3(n80), .A4(n44), .A5(n81), .A6(n65), 
        .Y(n93) );
  AO221X1_RVT U86 ( .A1(A[6]), .A2(n27), .A3(A[5]), .A4(n35), .A5(n94), .Y(n65) );
  AO22X1_RVT U87 ( .A1(A[8]), .A2(n34), .A3(A[7]), .A4(n30), .Y(n94) );
  AO221X1_RVT U88 ( .A1(A[10]), .A2(n27), .A3(A[9]), .A4(n36), .A5(n95), .Y(
        n44) );
  AO22X1_RVT U89 ( .A1(A[12]), .A2(n33), .A3(A[11]), .A4(n32), .Y(n95) );
  OA21X1_RVT U90 ( .A1(n96), .A2(n97), .A3(n75), .Y(n90) );
  AO22X1_RVT U91 ( .A1(A[1]), .A2(n36), .A3(A[2]), .A4(n28), .Y(n97) );
  AO22X1_RVT U92 ( .A1(A[4]), .A2(n34), .A3(A[3]), .A4(n32), .Y(n96) );
  AND2X1_RVT U93 ( .A1(n89), .A2(n77), .Y(B[19]) );
  AND2X1_RVT U94 ( .A1(n89), .A2(n85), .Y(B[18]) );
  AND2X1_RVT U95 ( .A1(n39), .A2(n98), .Y(n89) );
  AND2X1_RVT U96 ( .A1(n92), .A2(n98), .Y(B[17]) );
  AND2X1_RVT U97 ( .A1(n39), .A2(n46), .Y(n92) );
  MUX21X1_RVT U98 ( .A1(n68), .A2(n67), .S0(n40), .Y(n46) );
  AND2X1_RVT U99 ( .A1(n99), .A2(n98), .Y(B[16]) );
  AO222X1_RVT U100 ( .A1(n43), .A2(n57), .A3(n56), .A4(n35), .A5(n2), .A6(n25), 
        .Y(B[15]) );
  AO222X1_RVT U101 ( .A1(n63), .A2(n45), .A3(n43), .A4(n61), .A5(n2), .A6(n62), 
        .Y(B[14]) );
  AND2X1_RVT U102 ( .A1(n100), .A2(n40), .Y(n63) );
  AO222X1_RVT U103 ( .A1(n43), .A2(n47), .A3(n56), .A4(n68), .A5(n2), .A6(n67), 
        .Y(B[13]) );
  AO221X1_RVT U104 ( .A1(A[18]), .A2(n28), .A3(A[17]), .A4(n36), .A5(n101), 
        .Y(n67) );
  AO22X1_RVT U105 ( .A1(A[20]), .A2(n34), .A3(A[19]), .A4(n32), .Y(n101) );
  AO221X1_RVT U106 ( .A1(A[22]), .A2(n26), .A3(A[21]), .A4(n42), .A5(n31), .Y(
        n68) );
  AO221X1_RVT U107 ( .A1(A[14]), .A2(n28), .A3(A[13]), .A4(n36), .A5(n102), 
        .Y(n47) );
  AO22X1_RVT U108 ( .A1(A[16]), .A2(n34), .A3(A[15]), .A4(n31), .Y(n102) );
  AND2X1_RVT U109 ( .A1(n45), .A2(n40), .Y(n56) );
  AO222X1_RVT U110 ( .A1(n45), .A2(n77), .A3(n43), .A4(n52), .A5(n2), .A6(n57), 
        .Y(B[11]) );
  AO22X1_RVT U111 ( .A1(A[18]), .A2(n34), .A3(A[17]), .A4(n32), .Y(n103) );
  AO221X1_RVT U112 ( .A1(A[12]), .A2(n28), .A3(A[11]), .A4(n35), .A5(n104), 
        .Y(n52) );
  AO22X1_RVT U113 ( .A1(A[14]), .A2(n34), .A3(A[13]), .A4(n31), .Y(n104) );
  AO222X1_RVT U114 ( .A1(n45), .A2(n85), .A3(n43), .A4(n59), .A5(n2), .A6(n61), 
        .Y(B[10]) );
  AO221X1_RVT U115 ( .A1(A[15]), .A2(n27), .A3(A[14]), .A4(n35), .A5(n105), 
        .Y(n61) );
  AO22X1_RVT U116 ( .A1(A[17]), .A2(n34), .A3(A[16]), .A4(n30), .Y(n105) );
  AO221X1_RVT U117 ( .A1(A[11]), .A2(n26), .A3(A[10]), .A4(n35), .A5(n106), 
        .Y(n59) );
  AO22X1_RVT U118 ( .A1(A[13]), .A2(n34), .A3(A[12]), .A4(n30), .Y(n106) );
  MUX21X1_RVT U119 ( .A1(n100), .A2(n62), .S0(n40), .Y(n85) );
  AO221X1_RVT U120 ( .A1(A[19]), .A2(n26), .A3(n36), .A4(A[18]), .A5(n107), 
        .Y(n62) );
  AO22X1_RVT U121 ( .A1(n34), .A2(A[21]), .A3(A[20]), .A4(n32), .Y(n107) );
  AO21X1_RVT U122 ( .A1(A[22]), .A2(n41), .A3(n28), .Y(n100) );
  AND2X1_RVT U123 ( .A1(n98), .A2(n108), .Y(n45) );
  AND2X1_RVT U124 ( .A1(n38), .A2(n37), .Y(n98) );
  OA21X1_RVT U125 ( .A1(n109), .A2(n110), .A3(n37), .Y(B[0]) );
  MUX21X1_RVT U126 ( .A1(n99), .A2(n111), .S0(n38), .Y(n110) );
  AO222X1_RVT U127 ( .A1(n79), .A2(n50), .A3(n80), .A4(n48), .A5(n81), .A6(n69), .Y(n111) );
  AO221X1_RVT U128 ( .A1(A[5]), .A2(n27), .A3(A[4]), .A4(n35), .A5(n112), .Y(
        n69) );
  AO22X1_RVT U129 ( .A1(A[7]), .A2(n33), .A3(A[6]), .A4(n30), .Y(n112) );
  AND2X1_RVT U130 ( .A1(n39), .A2(SH[2]), .Y(n81) );
  AND2X1_RVT U131 ( .A1(n40), .A2(n108), .Y(n80) );
  AO221X1_RVT U132 ( .A1(A[13]), .A2(n26), .A3(A[12]), .A4(n35), .A5(n114), 
        .Y(n50) );
  AO22X1_RVT U133 ( .A1(A[15]), .A2(n34), .A3(A[14]), .A4(n30), .Y(n114) );
  AND2X1_RVT U134 ( .A1(SH[2]), .A2(n108), .Y(n79) );
  AND2X1_RVT U135 ( .A1(n39), .A2(n49), .Y(n99) );
  MUX21X1_RVT U136 ( .A1(n72), .A2(n71), .S0(n40), .Y(n49) );
  OA21X1_RVT U137 ( .A1(n115), .A2(n116), .A3(n75), .Y(n109) );
  AND3X1_RVT U138 ( .A1(n38), .A2(n40), .A3(n39), .Y(n75) );
  OR2X1_RVT U139 ( .A1(SH[3]), .A2(n117), .Y(n108) );
  OR2X1_RVT U140 ( .A1(SH[4]), .A2(n117), .Y(n88) );
  OR2X1_RVT U141 ( .A1(SH[5]), .A2(SH[6]), .Y(n117) );
  AO22X1_RVT U142 ( .A1(A[0]), .A2(n36), .A3(A[1]), .A4(n28), .Y(n116) );
  AO22X1_RVT U143 ( .A1(A[3]), .A2(n33), .A3(A[2]), .A4(n32), .Y(n115) );
endmodule


module FPU_CAL_DW01_sub_4 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [8:0] carry;

  FADDX1_RVT U2_7 ( .A(A[7]), .B(n1), .CI(carry[7]), .S(DIFF[7]) );
  FADDX1_RVT U2_6 ( .A(A[6]), .B(n2), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FADDX1_RVT U2_4 ( .A(A[4]), .B(n4), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FADDX1_RVT U2_3 ( .A(A[3]), .B(n5), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FADDX1_RVT U2_5 ( .A(A[5]), .B(n3), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FADDX1_RVT U2_2 ( .A(A[2]), .B(n6), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FADDX1_RVT U2_1 ( .A(A[1]), .B(n7), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  INVX1_RVT U1 ( .A(B[1]), .Y(n7) );
  INVX1_RVT U2 ( .A(B[0]), .Y(n8) );
  XNOR2X1_RVT U3 ( .A1(A[0]), .A2(n8), .Y(DIFF[0]) );
  OR2X1_RVT U4 ( .A1(n8), .A2(A[0]), .Y(carry[1]) );
  INVX1_RVT U5 ( .A(B[2]), .Y(n6) );
  INVX1_RVT U6 ( .A(B[5]), .Y(n3) );
  INVX1_RVT U7 ( .A(B[3]), .Y(n5) );
  INVX1_RVT U8 ( .A(B[4]), .Y(n4) );
  INVX1_RVT U9 ( .A(B[6]), .Y(n2) );
  INVX1_RVT U10 ( .A(B[7]), .Y(n1) );
endmodule


module FPU_CAL_DW_rash_1 ( A, DATA_TC, SH, SH_TC, B );
  input [23:0] A;
  input [7:0] SH;
  output [23:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116;

  INVX1_RVT U3 ( .A(SH[1]), .Y(n33) );
  INVX1_RVT U4 ( .A(SH[7]), .Y(n29) );
  INVX1_RVT U5 ( .A(n83), .Y(n30) );
  INVX1_RVT U6 ( .A(n17), .Y(n18) );
  INVX1_RVT U7 ( .A(n17), .Y(n19) );
  AND2X1_RVT U8 ( .A1(n74), .A2(n94), .Y(n1) );
  INVX1_RVT U9 ( .A(SH[2]), .Y(n32) );
  NAND2X0_RVT U10 ( .A1(n34), .A2(n33), .Y(n2) );
  NAND2X0_RVT U11 ( .A1(SH[0]), .A2(n33), .Y(n4) );
  AND2X1_RVT U12 ( .A1(n68), .A2(n29), .Y(n35) );
  INVX1_RVT U13 ( .A(n14), .Y(n15) );
  INVX1_RVT U14 ( .A(n22), .Y(n23) );
  INVX1_RVT U15 ( .A(n2), .Y(n27) );
  INVX1_RVT U16 ( .A(n2), .Y(n28) );
  INVX1_RVT U17 ( .A(n76), .Y(n24) );
  INVX1_RVT U18 ( .A(n76), .Y(n14) );
  INVX1_RVT U19 ( .A(n3), .Y(n26) );
  INVX1_RVT U20 ( .A(n4), .Y(n20) );
  AND2X1_RVT U21 ( .A1(n34), .A2(SH[1]), .Y(n22) );
  INVX1_RVT U22 ( .A(n3), .Y(n25) );
  AND2X1_RVT U23 ( .A1(n34), .A2(SH[1]), .Y(n76) );
  INVX1_RVT U24 ( .A(n4), .Y(n21) );
  NAND2X0_RVT U25 ( .A1(SH[0]), .A2(SH[1]), .Y(n3) );
  INVX1_RVT U26 ( .A(SH[0]), .Y(n34) );
  INVX1_RVT U27 ( .A(n14), .Y(n16) );
  INVX1_RVT U28 ( .A(n105), .Y(n31) );
  INVX1_RVT U29 ( .A(n24), .Y(n5) );
  NBUFFX2_RVT U30 ( .A(n5), .Y(n6) );
  NBUFFX2_RVT U31 ( .A(n5), .Y(n7) );
  NBUFFX2_RVT U32 ( .A(n5), .Y(n8) );
  NBUFFX2_RVT U33 ( .A(n5), .Y(n9) );
  NBUFFX2_RVT U34 ( .A(n5), .Y(n10) );
  INVX1_RVT U35 ( .A(n23), .Y(n11) );
  NBUFFX2_RVT U36 ( .A(n11), .Y(n12) );
  NBUFFX2_RVT U37 ( .A(n11), .Y(n13) );
  INVX1_RVT U38 ( .A(n22), .Y(n17) );
  AO222X1_RVT U39 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .A5(n1), .A6(n39), 
        .Y(B[9]) );
  AO222X1_RVT U40 ( .A1(n35), .A2(n40), .A3(n37), .A4(n41), .A5(n1), .A6(n42), 
        .Y(B[8]) );
  AO221X1_RVT U41 ( .A1(n35), .A2(n43), .A3(n1), .A4(n44), .A5(n45), .Y(B[7])
         );
  AO222X1_RVT U42 ( .A1(n46), .A2(n47), .A3(n48), .A4(n27), .A5(n49), .A6(n50), 
        .Y(n45) );
  AO221X1_RVT U43 ( .A1(n35), .A2(n51), .A3(n1), .A4(n52), .A5(n53), .Y(B[6])
         );
  AO222X1_RVT U44 ( .A1(n49), .A2(n54), .A3(n46), .A4(n55), .A5(n56), .A6(n57), 
        .Y(n53) );
  AO221X1_RVT U45 ( .A1(n35), .A2(n58), .A3(n1), .A4(n36), .A5(n59), .Y(B[5])
         );
  AO222X1_RVT U46 ( .A1(n46), .A2(n60), .A3(n48), .A4(n61), .A5(n49), .A6(n39), 
        .Y(n59) );
  AO221X1_RVT U47 ( .A1(n35), .A2(n62), .A3(n1), .A4(n40), .A5(n63), .Y(B[4])
         );
  AO222X1_RVT U48 ( .A1(n46), .A2(n64), .A3(n48), .A4(n65), .A5(n49), .A6(n42), 
        .Y(n63) );
  AND2X1_RVT U49 ( .A1(n57), .A2(n32), .Y(n48) );
  AND2X1_RVT U50 ( .A1(n66), .A2(n29), .Y(n57) );
  AND2X1_RVT U51 ( .A1(n37), .A2(SH[2]), .Y(n46) );
  AND2X1_RVT U52 ( .A1(n67), .A2(n29), .Y(B[3]) );
  AO222X1_RVT U53 ( .A1(n68), .A2(n69), .A3(n66), .A4(n70), .A5(n30), .A6(n71), 
        .Y(n67) );
  AO222X1_RVT U54 ( .A1(n72), .A2(n50), .A3(n73), .A4(n44), .A5(n74), .A6(n43), 
        .Y(n71) );
  AO221X1_RVT U55 ( .A1(A[8]), .A2(n21), .A3(A[7]), .A4(n27), .A5(n75), .Y(n43) );
  AO22X1_RVT U56 ( .A1(A[10]), .A2(n26), .A3(A[9]), .A4(n13), .Y(n75) );
  AO221X1_RVT U57 ( .A1(A[4]), .A2(n20), .A3(A[3]), .A4(n28), .A5(n77), .Y(n69) );
  AO22X1_RVT U58 ( .A1(A[6]), .A2(n25), .A3(A[5]), .A4(n16), .Y(n77) );
  AND2X1_RVT U59 ( .A1(n78), .A2(n29), .Y(B[2]) );
  AO222X1_RVT U60 ( .A1(n68), .A2(n79), .A3(n66), .A4(n80), .A5(n30), .A6(n81), 
        .Y(n78) );
  AO222X1_RVT U61 ( .A1(n72), .A2(n54), .A3(n73), .A4(n52), .A5(n74), .A6(n51), 
        .Y(n81) );
  AO221X1_RVT U62 ( .A1(A[7]), .A2(n21), .A3(A[6]), .A4(n28), .A5(n82), .Y(n51) );
  AO22X1_RVT U63 ( .A1(A[9]), .A2(n25), .A3(A[8]), .A4(n8), .Y(n82) );
  AND2X1_RVT U64 ( .A1(n31), .A2(n83), .Y(n66) );
  AO221X1_RVT U65 ( .A1(A[3]), .A2(n21), .A3(A[2]), .A4(n28), .A5(n84), .Y(n79) );
  AO22X1_RVT U66 ( .A1(A[5]), .A2(n26), .A3(A[4]), .A4(n9), .Y(n84) );
  AND2X1_RVT U67 ( .A1(n35), .A2(n28), .Y(B[23]) );
  AND2X1_RVT U68 ( .A1(n85), .A2(n56), .Y(B[22]) );
  AND2X1_RVT U69 ( .A1(n35), .A2(n61), .Y(B[21]) );
  AND2X1_RVT U70 ( .A1(n35), .A2(n65), .Y(B[20]) );
  OA21X1_RVT U71 ( .A1(n86), .A2(n87), .A3(n29), .Y(B[1]) );
  MUX21X1_RVT U72 ( .A1(n88), .A2(n89), .S0(n30), .Y(n87) );
  AO222X1_RVT U73 ( .A1(n72), .A2(n39), .A3(n73), .A4(n36), .A5(n74), .A6(n58), 
        .Y(n89) );
  AO221X1_RVT U74 ( .A1(A[6]), .A2(n21), .A3(A[5]), .A4(n27), .A5(n90), .Y(n58) );
  AO22X1_RVT U75 ( .A1(A[8]), .A2(n25), .A3(A[7]), .A4(n16), .Y(n90) );
  AO221X1_RVT U76 ( .A1(A[10]), .A2(n21), .A3(A[9]), .A4(n28), .A5(n91), .Y(
        n36) );
  AO22X1_RVT U77 ( .A1(A[12]), .A2(n25), .A3(A[11]), .A4(n7), .Y(n91) );
  OA21X1_RVT U78 ( .A1(n92), .A2(n93), .A3(n68), .Y(n86) );
  AO22X1_RVT U79 ( .A1(A[1]), .A2(n28), .A3(A[2]), .A4(n21), .Y(n93) );
  AO22X1_RVT U80 ( .A1(A[4]), .A2(n26), .A3(A[3]), .A4(n7), .Y(n92) );
  AND2X1_RVT U81 ( .A1(n85), .A2(n70), .Y(B[19]) );
  AND2X1_RVT U82 ( .A1(n85), .A2(n80), .Y(B[18]) );
  AND2X1_RVT U83 ( .A1(n31), .A2(n94), .Y(n85) );
  AND2X1_RVT U84 ( .A1(n88), .A2(n94), .Y(B[17]) );
  AND2X1_RVT U85 ( .A1(n31), .A2(n38), .Y(n88) );
  MUX21X1_RVT U86 ( .A1(n61), .A2(n60), .S0(n32), .Y(n38) );
  AND2X1_RVT U87 ( .A1(n95), .A2(n94), .Y(B[16]) );
  AO222X1_RVT U88 ( .A1(n35), .A2(n50), .A3(n49), .A4(n27), .A5(n1), .A6(n47), 
        .Y(B[15]) );
  AO222X1_RVT U89 ( .A1(n56), .A2(n37), .A3(n35), .A4(n54), .A5(n1), .A6(n55), 
        .Y(B[14]) );
  AND2X1_RVT U90 ( .A1(n96), .A2(n32), .Y(n56) );
  AO222X1_RVT U91 ( .A1(n35), .A2(n39), .A3(n49), .A4(n61), .A5(n1), .A6(n60), 
        .Y(B[13]) );
  AO221X1_RVT U92 ( .A1(A[18]), .A2(n21), .A3(A[17]), .A4(n28), .A5(n97), .Y(
        n60) );
  AO22X1_RVT U93 ( .A1(A[20]), .A2(n25), .A3(A[19]), .A4(n15), .Y(n97) );
  AO221X1_RVT U94 ( .A1(A[22]), .A2(n21), .A3(A[21]), .A4(n34), .A5(n16), .Y(
        n61) );
  AO221X1_RVT U95 ( .A1(A[14]), .A2(n21), .A3(A[13]), .A4(n28), .A5(n98), .Y(
        n39) );
  AO22X1_RVT U96 ( .A1(A[16]), .A2(n26), .A3(A[15]), .A4(n6), .Y(n98) );
  AO222X1_RVT U97 ( .A1(n35), .A2(n42), .A3(n49), .A4(n65), .A5(n1), .A6(n64), 
        .Y(B[12]) );
  AND2X1_RVT U98 ( .A1(n37), .A2(n32), .Y(n49) );
  AO222X1_RVT U99 ( .A1(n37), .A2(n70), .A3(n35), .A4(n44), .A5(n1), .A6(n50), 
        .Y(B[11]) );
  AO221X1_RVT U100 ( .A1(A[16]), .A2(n20), .A3(A[15]), .A4(n27), .A5(n99), .Y(
        n50) );
  AO22X1_RVT U101 ( .A1(A[18]), .A2(n26), .A3(A[17]), .A4(n15), .Y(n99) );
  AO221X1_RVT U102 ( .A1(A[12]), .A2(n20), .A3(A[11]), .A4(n27), .A5(n100), 
        .Y(n44) );
  AO22X1_RVT U103 ( .A1(A[14]), .A2(n25), .A3(A[13]), .A4(n12), .Y(n100) );
  MUX21X1_RVT U104 ( .A1(n28), .A2(n47), .S0(n32), .Y(n70) );
  AO221X1_RVT U105 ( .A1(A[20]), .A2(n21), .A3(n28), .A4(A[19]), .A5(n101), 
        .Y(n47) );
  AO22X1_RVT U106 ( .A1(n26), .A2(A[22]), .A3(n10), .A4(A[21]), .Y(n101) );
  AO222X1_RVT U107 ( .A1(n37), .A2(n80), .A3(n35), .A4(n52), .A5(n1), .A6(n54), 
        .Y(B[10]) );
  AO221X1_RVT U108 ( .A1(A[15]), .A2(n21), .A3(A[14]), .A4(n27), .A5(n102), 
        .Y(n54) );
  AO22X1_RVT U109 ( .A1(A[17]), .A2(n26), .A3(A[16]), .A4(n8), .Y(n102) );
  AO221X1_RVT U110 ( .A1(A[11]), .A2(n20), .A3(A[10]), .A4(n27), .A5(n103), 
        .Y(n52) );
  AO22X1_RVT U111 ( .A1(A[13]), .A2(n26), .A3(A[12]), .A4(n9), .Y(n103) );
  MUX21X1_RVT U112 ( .A1(n96), .A2(n55), .S0(n32), .Y(n80) );
  AO221X1_RVT U113 ( .A1(A[19]), .A2(n20), .A3(n28), .A4(A[18]), .A5(n104), 
        .Y(n55) );
  AO22X1_RVT U114 ( .A1(n25), .A2(A[21]), .A3(A[20]), .A4(n6), .Y(n104) );
  AO21X1_RVT U115 ( .A1(A[22]), .A2(n33), .A3(n20), .Y(n96) );
  AND2X1_RVT U116 ( .A1(n94), .A2(n105), .Y(n37) );
  AND2X1_RVT U117 ( .A1(n30), .A2(n29), .Y(n94) );
  OA21X1_RVT U118 ( .A1(n106), .A2(n107), .A3(n29), .Y(B[0]) );
  MUX21X1_RVT U119 ( .A1(n95), .A2(n108), .S0(n30), .Y(n107) );
  AO222X1_RVT U120 ( .A1(n72), .A2(n42), .A3(n73), .A4(n40), .A5(n74), .A6(n62), .Y(n108) );
  AO221X1_RVT U121 ( .A1(A[5]), .A2(n20), .A3(A[4]), .A4(n27), .A5(n109), .Y(
        n62) );
  AO22X1_RVT U122 ( .A1(A[7]), .A2(n25), .A3(A[6]), .A4(n15), .Y(n109) );
  AND2X1_RVT U123 ( .A1(n31), .A2(SH[2]), .Y(n74) );
  AO221X1_RVT U124 ( .A1(A[9]), .A2(n21), .A3(A[8]), .A4(n27), .A5(n110), .Y(
        n40) );
  AO22X1_RVT U125 ( .A1(A[11]), .A2(n25), .A3(A[10]), .A4(n11), .Y(n110) );
  AND2X1_RVT U126 ( .A1(n32), .A2(n105), .Y(n73) );
  AO221X1_RVT U127 ( .A1(A[13]), .A2(n20), .A3(A[12]), .A4(n27), .A5(n111), 
        .Y(n42) );
  AO22X1_RVT U128 ( .A1(A[15]), .A2(n26), .A3(A[14]), .A4(n18), .Y(n111) );
  AND2X1_RVT U129 ( .A1(SH[2]), .A2(n105), .Y(n72) );
  AND2X1_RVT U130 ( .A1(n31), .A2(n41), .Y(n95) );
  MUX21X1_RVT U131 ( .A1(n65), .A2(n64), .S0(n32), .Y(n41) );
  AO221X1_RVT U132 ( .A1(A[17]), .A2(n20), .A3(A[16]), .A4(n27), .A5(n112), 
        .Y(n64) );
  AO22X1_RVT U133 ( .A1(n25), .A2(A[19]), .A3(A[18]), .A4(n19), .Y(n112) );
  AO221X1_RVT U134 ( .A1(A[21]), .A2(SH[0]), .A3(A[22]), .A4(SH[1]), .A5(n113), 
        .Y(n65) );
  AO21X1_RVT U135 ( .A1(n28), .A2(A[20]), .A3(n25), .Y(n113) );
  OA21X1_RVT U136 ( .A1(n114), .A2(n115), .A3(n68), .Y(n106) );
  AND3X1_RVT U137 ( .A1(n30), .A2(n32), .A3(n31), .Y(n68) );
  OR2X1_RVT U138 ( .A1(SH[3]), .A2(n116), .Y(n105) );
  OR2X1_RVT U139 ( .A1(SH[4]), .A2(n116), .Y(n83) );
  OR2X1_RVT U140 ( .A1(SH[5]), .A2(SH[6]), .Y(n116) );
  AO22X1_RVT U141 ( .A1(A[0]), .A2(n28), .A3(A[1]), .A4(n21), .Y(n115) );
  AO22X1_RVT U142 ( .A1(A[3]), .A2(n25), .A3(A[2]), .A4(n10), .Y(n114) );
endmodule


module FPU_CAL_DW01_sub_5 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [8:0] carry;

  FADDX1_RVT U2_1 ( .A(A[1]), .B(n7), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  FADDX1_RVT U2_4 ( .A(A[4]), .B(n4), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FADDX1_RVT U2_5 ( .A(A[5]), .B(n3), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FADDX1_RVT U2_2 ( .A(A[2]), .B(n6), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FADDX1_RVT U2_3 ( .A(A[3]), .B(n5), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FADDX1_RVT U2_7 ( .A(A[7]), .B(n1), .CI(carry[7]), .S(DIFF[7]) );
  FADDX1_RVT U2_6 ( .A(A[6]), .B(n2), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FADDX1_RVT U2_0 ( .A(A[0]), .B(n8), .CI(1'b1), .CO(carry[1]), .S(DIFF[0]) );
  INVX1_RVT U1 ( .A(B[0]), .Y(n8) );
  INVX1_RVT U2 ( .A(B[1]), .Y(n7) );
  INVX1_RVT U3 ( .A(B[3]), .Y(n5) );
  INVX1_RVT U4 ( .A(B[5]), .Y(n3) );
  INVX1_RVT U5 ( .A(B[2]), .Y(n6) );
  INVX1_RVT U6 ( .A(B[4]), .Y(n4) );
  INVX1_RVT U7 ( .A(B[6]), .Y(n2) );
  INVX1_RVT U8 ( .A(B[7]), .Y(n1) );
endmodule


module FPU_CAL_DW01_add_4 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  AND2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
  XOR2X1_RVT U2 ( .A1(B[8]), .A2(carry[8]), .Y(SUM[8]) );
  XOR2X1_RVT U3 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
endmodule


module FPU_CAL_DW01_add_2 ( A, B, CI, SUM, CO );
  input [45:0] A;
  input [45:0] B;
  output [45:0] SUM;
  input CI;
  output CO;
  wire   \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , \A[17] , \A[16] ,
         \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] ,
         \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110;
  assign SUM[22] = \A[22] ;
  assign \A[22]  = A[22];
  assign SUM[21] = \A[21] ;
  assign \A[21]  = A[21];
  assign SUM[20] = \A[20] ;
  assign \A[20]  = A[20];
  assign SUM[19] = \A[19] ;
  assign \A[19]  = A[19];
  assign SUM[18] = \A[18] ;
  assign \A[18]  = A[18];
  assign SUM[17] = \A[17] ;
  assign \A[17]  = A[17];
  assign SUM[16] = \A[16] ;
  assign \A[16]  = A[16];
  assign SUM[15] = \A[15] ;
  assign \A[15]  = A[15];
  assign SUM[14] = \A[14] ;
  assign \A[14]  = A[14];
  assign SUM[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign SUM[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign SUM[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign SUM[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  INVX1_RVT U2 ( .A(n109), .Y(n24) );
  INVX1_RVT U3 ( .A(n94), .Y(n19) );
  INVX1_RVT U4 ( .A(n97), .Y(n20) );
  INVX1_RVT U5 ( .A(n104), .Y(n22) );
  INVX1_RVT U6 ( .A(n107), .Y(n23) );
  INVX1_RVT U7 ( .A(n90), .Y(n18) );
  INVX1_RVT U8 ( .A(n86), .Y(n17) );
  INVX1_RVT U9 ( .A(n30), .Y(n3) );
  INVX1_RVT U10 ( .A(n38), .Y(n5) );
  INVX1_RVT U11 ( .A(n70), .Y(n13) );
  INVX1_RVT U12 ( .A(n54), .Y(n9) );
  INVX1_RVT U13 ( .A(n74), .Y(n14) );
  INVX1_RVT U14 ( .A(n42), .Y(n6) );
  INVX1_RVT U15 ( .A(n78), .Y(n15) );
  INVX1_RVT U16 ( .A(n62), .Y(n11) );
  INVX1_RVT U17 ( .A(n58), .Y(n10) );
  INVX1_RVT U18 ( .A(n46), .Y(n7) );
  INVX1_RVT U19 ( .A(n82), .Y(n16) );
  INVX1_RVT U20 ( .A(n34), .Y(n4) );
  INVX1_RVT U21 ( .A(n66), .Y(n12) );
  INVX1_RVT U22 ( .A(n50), .Y(n8) );
  INVX1_RVT U23 ( .A(n96), .Y(n21) );
  XNOR2X1_RVT U24 ( .A1(B[45]), .A2(n25), .Y(SUM[45]) );
  INVX1_RVT U25 ( .A(B[44]), .Y(n2) );
  AND2X1_RVT U26 ( .A1(n110), .A2(n109), .Y(SUM[23]) );
  OA22X1_RVT U27 ( .A1(n26), .A2(n2), .A3(n27), .A4(B[45]), .Y(n25) );
  AND2X1_RVT U28 ( .A1(n27), .A2(B[45]), .Y(n26) );
  XNOR3X1_RVT U29 ( .A1(B[44]), .A2(A[44]), .A3(n27), .Y(SUM[44]) );
  OA21X1_RVT U30 ( .A1(n28), .A2(n3), .A3(n29), .Y(n27) );
  XOR2X1_RVT U31 ( .A1(n31), .A2(n28), .Y(SUM[43]) );
  OA21X1_RVT U32 ( .A1(n32), .A2(n4), .A3(n33), .Y(n28) );
  NAND2X0_RVT U33 ( .A1(n30), .A2(n29), .Y(n31) );
  NAND2X0_RVT U34 ( .A1(B[43]), .A2(A[43]), .Y(n29) );
  OR2X1_RVT U35 ( .A1(B[43]), .A2(A[43]), .Y(n30) );
  XOR2X1_RVT U36 ( .A1(n35), .A2(n32), .Y(SUM[42]) );
  OA21X1_RVT U37 ( .A1(n36), .A2(n5), .A3(n37), .Y(n32) );
  NAND2X0_RVT U38 ( .A1(n34), .A2(n33), .Y(n35) );
  NAND2X0_RVT U39 ( .A1(B[42]), .A2(A[42]), .Y(n33) );
  OR2X1_RVT U40 ( .A1(B[42]), .A2(A[42]), .Y(n34) );
  XOR2X1_RVT U41 ( .A1(n39), .A2(n36), .Y(SUM[41]) );
  OA21X1_RVT U42 ( .A1(n40), .A2(n6), .A3(n41), .Y(n36) );
  NAND2X0_RVT U43 ( .A1(n38), .A2(n37), .Y(n39) );
  NAND2X0_RVT U44 ( .A1(B[41]), .A2(A[41]), .Y(n37) );
  OR2X1_RVT U45 ( .A1(B[41]), .A2(A[41]), .Y(n38) );
  XOR2X1_RVT U46 ( .A1(n43), .A2(n40), .Y(SUM[40]) );
  OA21X1_RVT U47 ( .A1(n44), .A2(n7), .A3(n45), .Y(n40) );
  NAND2X0_RVT U48 ( .A1(n42), .A2(n41), .Y(n43) );
  NAND2X0_RVT U49 ( .A1(B[40]), .A2(A[40]), .Y(n41) );
  OR2X1_RVT U50 ( .A1(B[40]), .A2(A[40]), .Y(n42) );
  XOR2X1_RVT U51 ( .A1(n47), .A2(n44), .Y(SUM[39]) );
  OA21X1_RVT U52 ( .A1(n48), .A2(n8), .A3(n49), .Y(n44) );
  NAND2X0_RVT U53 ( .A1(n46), .A2(n45), .Y(n47) );
  NAND2X0_RVT U54 ( .A1(B[39]), .A2(A[39]), .Y(n45) );
  OR2X1_RVT U55 ( .A1(B[39]), .A2(A[39]), .Y(n46) );
  XOR2X1_RVT U56 ( .A1(n51), .A2(n48), .Y(SUM[38]) );
  OA21X1_RVT U57 ( .A1(n52), .A2(n9), .A3(n53), .Y(n48) );
  NAND2X0_RVT U58 ( .A1(n50), .A2(n49), .Y(n51) );
  NAND2X0_RVT U59 ( .A1(B[38]), .A2(A[38]), .Y(n49) );
  OR2X1_RVT U60 ( .A1(B[38]), .A2(A[38]), .Y(n50) );
  XOR2X1_RVT U61 ( .A1(n55), .A2(n52), .Y(SUM[37]) );
  OA21X1_RVT U62 ( .A1(n56), .A2(n10), .A3(n57), .Y(n52) );
  NAND2X0_RVT U63 ( .A1(n54), .A2(n53), .Y(n55) );
  NAND2X0_RVT U64 ( .A1(B[37]), .A2(A[37]), .Y(n53) );
  OR2X1_RVT U65 ( .A1(B[37]), .A2(A[37]), .Y(n54) );
  XOR2X1_RVT U66 ( .A1(n59), .A2(n56), .Y(SUM[36]) );
  OA21X1_RVT U67 ( .A1(n60), .A2(n11), .A3(n61), .Y(n56) );
  NAND2X0_RVT U68 ( .A1(n58), .A2(n57), .Y(n59) );
  NAND2X0_RVT U69 ( .A1(B[36]), .A2(A[36]), .Y(n57) );
  OR2X1_RVT U70 ( .A1(B[36]), .A2(A[36]), .Y(n58) );
  XOR2X1_RVT U71 ( .A1(n63), .A2(n60), .Y(SUM[35]) );
  OA21X1_RVT U72 ( .A1(n64), .A2(n12), .A3(n65), .Y(n60) );
  NAND2X0_RVT U73 ( .A1(n62), .A2(n61), .Y(n63) );
  NAND2X0_RVT U74 ( .A1(B[35]), .A2(A[35]), .Y(n61) );
  OR2X1_RVT U75 ( .A1(B[35]), .A2(A[35]), .Y(n62) );
  XOR2X1_RVT U76 ( .A1(n67), .A2(n64), .Y(SUM[34]) );
  OA21X1_RVT U77 ( .A1(n68), .A2(n13), .A3(n69), .Y(n64) );
  NAND2X0_RVT U78 ( .A1(n66), .A2(n65), .Y(n67) );
  NAND2X0_RVT U79 ( .A1(B[34]), .A2(A[34]), .Y(n65) );
  OR2X1_RVT U80 ( .A1(B[34]), .A2(A[34]), .Y(n66) );
  XOR2X1_RVT U81 ( .A1(n71), .A2(n68), .Y(SUM[33]) );
  OA21X1_RVT U82 ( .A1(n72), .A2(n14), .A3(n73), .Y(n68) );
  NAND2X0_RVT U83 ( .A1(n70), .A2(n69), .Y(n71) );
  NAND2X0_RVT U84 ( .A1(B[33]), .A2(A[33]), .Y(n69) );
  OR2X1_RVT U85 ( .A1(B[33]), .A2(A[33]), .Y(n70) );
  XOR2X1_RVT U86 ( .A1(n75), .A2(n72), .Y(SUM[32]) );
  OA21X1_RVT U87 ( .A1(n76), .A2(n15), .A3(n77), .Y(n72) );
  NAND2X0_RVT U88 ( .A1(n74), .A2(n73), .Y(n75) );
  NAND2X0_RVT U89 ( .A1(B[32]), .A2(A[32]), .Y(n73) );
  OR2X1_RVT U90 ( .A1(B[32]), .A2(A[32]), .Y(n74) );
  XOR2X1_RVT U91 ( .A1(n79), .A2(n76), .Y(SUM[31]) );
  OA21X1_RVT U92 ( .A1(n80), .A2(n16), .A3(n81), .Y(n76) );
  NAND2X0_RVT U93 ( .A1(n78), .A2(n77), .Y(n79) );
  NAND2X0_RVT U94 ( .A1(B[31]), .A2(A[31]), .Y(n77) );
  OR2X1_RVT U95 ( .A1(B[31]), .A2(A[31]), .Y(n78) );
  XOR2X1_RVT U96 ( .A1(n83), .A2(n80), .Y(SUM[30]) );
  OA21X1_RVT U97 ( .A1(n84), .A2(n17), .A3(n85), .Y(n80) );
  NAND2X0_RVT U98 ( .A1(n82), .A2(n81), .Y(n83) );
  NAND2X0_RVT U99 ( .A1(B[30]), .A2(A[30]), .Y(n81) );
  OR2X1_RVT U100 ( .A1(B[30]), .A2(A[30]), .Y(n82) );
  XOR2X1_RVT U101 ( .A1(n87), .A2(n84), .Y(SUM[29]) );
  AOI21X1_RVT U102 ( .A1(n88), .A2(n89), .A3(n18), .Y(n84) );
  NAND2X0_RVT U103 ( .A1(n86), .A2(n85), .Y(n87) );
  NAND2X0_RVT U104 ( .A1(B[29]), .A2(A[29]), .Y(n85) );
  OR2X1_RVT U105 ( .A1(B[29]), .A2(A[29]), .Y(n86) );
  XNOR2X1_RVT U106 ( .A1(n91), .A2(n88), .Y(SUM[28]) );
  AO21X1_RVT U107 ( .A1(n92), .A2(n93), .A3(n19), .Y(n88) );
  AO21X1_RVT U108 ( .A1(n95), .A2(n96), .A3(n20), .Y(n92) );
  AO21X1_RVT U109 ( .A1(n98), .A2(n99), .A3(n22), .Y(n95) );
  NAND2X0_RVT U110 ( .A1(n89), .A2(n90), .Y(n91) );
  NAND2X0_RVT U111 ( .A1(B[28]), .A2(A[28]), .Y(n90) );
  OR2X1_RVT U112 ( .A1(B[28]), .A2(A[28]), .Y(n89) );
  XOR2X1_RVT U113 ( .A1(n100), .A2(n101), .Y(SUM[27]) );
  OA21X1_RVT U114 ( .A1(n21), .A2(n102), .A3(n97), .Y(n101) );
  NAND2X0_RVT U115 ( .A1(n93), .A2(n94), .Y(n100) );
  NAND2X0_RVT U116 ( .A1(B[27]), .A2(A[27]), .Y(n94) );
  OR2X1_RVT U117 ( .A1(B[27]), .A2(A[27]), .Y(n93) );
  XOR2X1_RVT U118 ( .A1(n103), .A2(n102), .Y(SUM[26]) );
  AOI21X1_RVT U119 ( .A1(n98), .A2(n99), .A3(n22), .Y(n102) );
  NAND2X0_RVT U120 ( .A1(n96), .A2(n97), .Y(n103) );
  NAND2X0_RVT U121 ( .A1(B[26]), .A2(A[26]), .Y(n97) );
  OR2X1_RVT U122 ( .A1(B[26]), .A2(A[26]), .Y(n96) );
  XNOR2X1_RVT U123 ( .A1(n105), .A2(n98), .Y(SUM[25]) );
  AO21X1_RVT U124 ( .A1(n24), .A2(n106), .A3(n23), .Y(n98) );
  NAND2X0_RVT U125 ( .A1(n99), .A2(n104), .Y(n105) );
  NAND2X0_RVT U126 ( .A1(B[25]), .A2(A[25]), .Y(n104) );
  OR2X1_RVT U127 ( .A1(B[25]), .A2(A[25]), .Y(n99) );
  XNOR2X1_RVT U128 ( .A1(n108), .A2(n24), .Y(SUM[24]) );
  NAND2X0_RVT U129 ( .A1(n106), .A2(n107), .Y(n108) );
  NAND2X0_RVT U130 ( .A1(B[24]), .A2(A[24]), .Y(n107) );
  OR2X1_RVT U131 ( .A1(B[24]), .A2(A[24]), .Y(n106) );
  NAND2X0_RVT U132 ( .A1(B[23]), .A2(A[23]), .Y(n109) );
  OR2X1_RVT U133 ( .A1(B[23]), .A2(A[23]), .Y(n110) );
endmodule


module FPU_CAL_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [23:0] A;
  input [23:0] B;
  output [47:0] PRODUCT;
  input TC;
  wire   \ab[23][22] , \ab[23][21] , \ab[23][20] , \ab[23][19] , \ab[23][18] ,
         \ab[23][17] , \ab[23][16] , \ab[23][15] , \ab[23][14] , \ab[23][13] ,
         \ab[23][12] , \ab[23][11] , \ab[23][10] , \ab[23][9] , \ab[23][8] ,
         \ab[23][7] , \ab[23][6] , \ab[23][5] , \ab[23][4] , \ab[23][3] ,
         \ab[23][2] , \ab[23][1] , \ab[23][0] , \ab[22][23] , \ab[22][22] ,
         \ab[22][21] , \ab[22][20] , \ab[22][19] , \ab[22][18] , \ab[22][17] ,
         \ab[22][16] , \ab[22][15] , \ab[22][14] , \ab[22][13] , \ab[22][12] ,
         \ab[22][11] , \ab[22][10] , \ab[22][9] , \ab[22][8] , \ab[22][7] ,
         \ab[22][6] , \ab[22][5] , \ab[22][4] , \ab[22][3] , \ab[22][2] ,
         \ab[22][1] , \ab[22][0] , \ab[21][23] , \ab[21][22] , \ab[21][21] ,
         \ab[21][20] , \ab[21][19] , \ab[21][18] , \ab[21][17] , \ab[21][16] ,
         \ab[21][15] , \ab[21][14] , \ab[21][13] , \ab[21][12] , \ab[21][11] ,
         \ab[21][10] , \ab[21][9] , \ab[21][8] , \ab[21][7] , \ab[21][6] ,
         \ab[21][5] , \ab[21][4] , \ab[21][3] , \ab[21][2] , \ab[21][1] ,
         \ab[21][0] , \ab[20][23] , \ab[20][22] , \ab[20][21] , \ab[20][20] ,
         \ab[20][19] , \ab[20][18] , \ab[20][17] , \ab[20][16] , \ab[20][15] ,
         \ab[20][14] , \ab[20][13] , \ab[20][12] , \ab[20][11] , \ab[20][10] ,
         \ab[20][9] , \ab[20][8] , \ab[20][7] , \ab[20][6] , \ab[20][5] ,
         \ab[20][4] , \ab[20][3] , \ab[20][2] , \ab[20][1] , \ab[20][0] ,
         \ab[19][23] , \ab[19][22] , \ab[19][21] , \ab[19][20] , \ab[19][19] ,
         \ab[19][18] , \ab[19][17] , \ab[19][16] , \ab[19][15] , \ab[19][14] ,
         \ab[19][13] , \ab[19][12] , \ab[19][11] , \ab[19][10] , \ab[19][9] ,
         \ab[19][8] , \ab[19][7] , \ab[19][6] , \ab[19][5] , \ab[19][4] ,
         \ab[19][3] , \ab[19][2] , \ab[19][1] , \ab[19][0] , \ab[18][23] ,
         \ab[18][22] , \ab[18][21] , \ab[18][20] , \ab[18][19] , \ab[18][18] ,
         \ab[18][17] , \ab[18][16] , \ab[18][15] , \ab[18][14] , \ab[18][13] ,
         \ab[18][12] , \ab[18][11] , \ab[18][10] , \ab[18][9] , \ab[18][8] ,
         \ab[18][7] , \ab[18][6] , \ab[18][5] , \ab[18][4] , \ab[18][3] ,
         \ab[18][2] , \ab[18][1] , \ab[18][0] , \ab[17][23] , \ab[17][22] ,
         \ab[17][21] , \ab[17][20] , \ab[17][19] , \ab[17][18] , \ab[17][17] ,
         \ab[17][16] , \ab[17][15] , \ab[17][14] , \ab[17][13] , \ab[17][12] ,
         \ab[17][11] , \ab[17][10] , \ab[17][9] , \ab[17][8] , \ab[17][7] ,
         \ab[17][6] , \ab[17][5] , \ab[17][4] , \ab[17][3] , \ab[17][2] ,
         \ab[17][1] , \ab[17][0] , \ab[16][23] , \ab[16][22] , \ab[16][21] ,
         \ab[16][20] , \ab[16][19] , \ab[16][18] , \ab[16][17] , \ab[16][16] ,
         \ab[16][15] , \ab[16][14] , \ab[16][13] , \ab[16][12] , \ab[16][11] ,
         \ab[16][10] , \ab[16][9] , \ab[16][8] , \ab[16][7] , \ab[16][6] ,
         \ab[16][5] , \ab[16][4] , \ab[16][3] , \ab[16][2] , \ab[16][1] ,
         \ab[16][0] , \ab[15][23] , \ab[15][22] , \ab[15][21] , \ab[15][20] ,
         \ab[15][19] , \ab[15][18] , \ab[15][17] , \ab[15][16] , \ab[15][15] ,
         \ab[15][14] , \ab[15][13] , \ab[15][12] , \ab[15][11] , \ab[15][10] ,
         \ab[15][9] , \ab[15][8] , \ab[15][7] , \ab[15][6] , \ab[15][5] ,
         \ab[15][4] , \ab[15][3] , \ab[15][2] , \ab[15][1] , \ab[15][0] ,
         \ab[14][23] , \ab[14][22] , \ab[14][21] , \ab[14][20] , \ab[14][19] ,
         \ab[14][18] , \ab[14][17] , \ab[14][16] , \ab[14][15] , \ab[14][14] ,
         \ab[14][13] , \ab[14][12] , \ab[14][11] , \ab[14][10] , \ab[14][9] ,
         \ab[14][8] , \ab[14][7] , \ab[14][6] , \ab[14][5] , \ab[14][4] ,
         \ab[14][3] , \ab[14][2] , \ab[14][1] , \ab[14][0] , \ab[13][23] ,
         \ab[13][22] , \ab[13][21] , \ab[13][20] , \ab[13][19] , \ab[13][18] ,
         \ab[13][17] , \ab[13][16] , \ab[13][15] , \ab[13][14] , \ab[13][13] ,
         \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] , \ab[13][8] ,
         \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] , \ab[13][3] ,
         \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][23] , \ab[12][22] ,
         \ab[12][21] , \ab[12][20] , \ab[12][19] , \ab[12][18] , \ab[12][17] ,
         \ab[12][16] , \ab[12][15] , \ab[12][14] , \ab[12][13] , \ab[12][12] ,
         \ab[12][11] , \ab[12][10] , \ab[12][9] , \ab[12][8] , \ab[12][7] ,
         \ab[12][6] , \ab[12][5] , \ab[12][4] , \ab[12][3] , \ab[12][2] ,
         \ab[12][1] , \ab[12][0] , \ab[11][23] , \ab[11][22] , \ab[11][21] ,
         \ab[11][20] , \ab[11][19] , \ab[11][18] , \ab[11][17] , \ab[11][16] ,
         \ab[11][15] , \ab[11][14] , \ab[11][13] , \ab[11][12] , \ab[11][11] ,
         \ab[11][10] , \ab[11][9] , \ab[11][8] , \ab[11][7] , \ab[11][6] ,
         \ab[11][5] , \ab[11][4] , \ab[11][3] , \ab[11][2] , \ab[11][1] ,
         \ab[11][0] , \ab[10][23] , \ab[10][22] , \ab[10][21] , \ab[10][20] ,
         \ab[10][19] , \ab[10][18] , \ab[10][17] , \ab[10][16] , \ab[10][15] ,
         \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] , \ab[10][10] ,
         \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] , \ab[10][5] ,
         \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] , \ab[10][0] ,
         \ab[9][23] , \ab[9][22] , \ab[9][21] , \ab[9][20] , \ab[9][19] ,
         \ab[9][18] , \ab[9][17] , \ab[9][16] , \ab[9][15] , \ab[9][14] ,
         \ab[9][13] , \ab[9][12] , \ab[9][11] , \ab[9][10] , \ab[9][9] ,
         \ab[9][8] , \ab[9][7] , \ab[9][6] , \ab[9][5] , \ab[9][4] ,
         \ab[9][3] , \ab[9][2] , \ab[9][1] , \ab[9][0] , \ab[8][23] ,
         \ab[8][22] , \ab[8][21] , \ab[8][20] , \ab[8][19] , \ab[8][18] ,
         \ab[8][17] , \ab[8][16] , \ab[8][15] , \ab[8][14] , \ab[8][13] ,
         \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] , \ab[8][8] ,
         \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] ,
         \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][23] , \ab[7][22] ,
         \ab[7][21] , \ab[7][20] , \ab[7][19] , \ab[7][18] , \ab[7][17] ,
         \ab[7][16] , \ab[7][15] , \ab[7][14] , \ab[7][13] , \ab[7][12] ,
         \ab[7][11] , \ab[7][10] , \ab[7][9] , \ab[7][8] , \ab[7][7] ,
         \ab[7][6] , \ab[7][5] , \ab[7][4] , \ab[7][3] , \ab[7][2] ,
         \ab[7][1] , \ab[7][0] , \ab[6][23] , \ab[6][22] , \ab[6][21] ,
         \ab[6][20] , \ab[6][19] , \ab[6][18] , \ab[6][17] , \ab[6][16] ,
         \ab[6][15] , \ab[6][14] , \ab[6][13] , \ab[6][12] , \ab[6][11] ,
         \ab[6][10] , \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] ,
         \ab[6][5] , \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] ,
         \ab[6][0] , \ab[5][23] , \ab[5][22] , \ab[5][21] , \ab[5][20] ,
         \ab[5][19] , \ab[5][18] , \ab[5][17] , \ab[5][16] , \ab[5][15] ,
         \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] , \ab[5][10] ,
         \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] , \ab[5][5] ,
         \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] , \ab[5][0] ,
         \ab[4][23] , \ab[4][22] , \ab[4][21] , \ab[4][20] , \ab[4][19] ,
         \ab[4][18] , \ab[4][17] , \ab[4][16] , \ab[4][15] , \ab[4][14] ,
         \ab[4][13] , \ab[4][12] , \ab[4][11] , \ab[4][10] , \ab[4][9] ,
         \ab[4][8] , \ab[4][7] , \ab[4][6] , \ab[4][5] , \ab[4][4] ,
         \ab[4][3] , \ab[4][2] , \ab[4][1] , \ab[4][0] , \ab[3][23] ,
         \ab[3][22] , \ab[3][21] , \ab[3][20] , \ab[3][19] , \ab[3][18] ,
         \ab[3][17] , \ab[3][16] , \ab[3][15] , \ab[3][14] , \ab[3][13] ,
         \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] , \ab[3][8] ,
         \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][23] , \ab[2][22] ,
         \ab[2][21] , \ab[2][20] , \ab[2][19] , \ab[2][18] , \ab[2][17] ,
         \ab[2][16] , \ab[2][15] , \ab[2][14] , \ab[2][13] , \ab[2][12] ,
         \ab[2][11] , \ab[2][10] , \ab[2][9] , \ab[2][8] , \ab[2][7] ,
         \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] , \ab[2][2] ,
         \ab[2][1] , \ab[2][0] , \ab[1][23] , \ab[1][22] , \ab[1][21] ,
         \ab[1][20] , \ab[1][19] , \ab[1][18] , \ab[1][17] , \ab[1][16] ,
         \ab[1][15] , \ab[1][14] , \ab[1][13] , \ab[1][12] , \ab[1][11] ,
         \ab[1][10] , \ab[1][9] , \ab[1][8] , \ab[1][7] , \ab[1][6] ,
         \ab[1][5] , \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] ,
         \ab[1][0] , \ab[0][23] , \ab[0][22] , \ab[0][21] , \ab[0][20] ,
         \ab[0][19] , \ab[0][18] , \ab[0][17] , \ab[0][16] , \ab[0][15] ,
         \ab[0][14] , \ab[0][13] , \ab[0][12] , \ab[0][11] , \ab[0][10] ,
         \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] ,
         \ab[0][4] , \ab[0][3] , \ab[0][2] , \ab[0][1] , \CARRYB[23][22] ,
         \CARRYB[23][21] , \CARRYB[23][20] , \CARRYB[23][19] ,
         \CARRYB[23][18] , \CARRYB[23][17] , \CARRYB[23][16] ,
         \CARRYB[23][15] , \CARRYB[23][14] , \CARRYB[23][13] ,
         \CARRYB[23][12] , \CARRYB[23][11] , \CARRYB[23][10] , \CARRYB[23][9] ,
         \CARRYB[23][8] , \CARRYB[23][7] , \CARRYB[23][6] , \CARRYB[23][5] ,
         \CARRYB[23][4] , \CARRYB[23][3] , \CARRYB[23][2] , \CARRYB[23][1] ,
         \CARRYB[23][0] , \CARRYB[22][22] , \CARRYB[22][21] , \CARRYB[22][20] ,
         \CARRYB[22][19] , \CARRYB[22][18] , \CARRYB[22][17] ,
         \CARRYB[22][16] , \CARRYB[22][15] , \CARRYB[22][14] ,
         \CARRYB[22][13] , \CARRYB[22][12] , \CARRYB[22][11] ,
         \CARRYB[22][10] , \CARRYB[22][9] , \CARRYB[22][8] , \CARRYB[22][7] ,
         \CARRYB[22][6] , \CARRYB[22][5] , \CARRYB[22][4] , \CARRYB[22][3] ,
         \CARRYB[22][2] , \CARRYB[22][1] , \CARRYB[22][0] , \CARRYB[21][22] ,
         \CARRYB[21][21] , \CARRYB[21][20] , \CARRYB[21][19] ,
         \CARRYB[21][18] , \CARRYB[21][17] , \CARRYB[21][16] ,
         \CARRYB[21][15] , \CARRYB[21][14] , \CARRYB[21][13] ,
         \CARRYB[21][12] , \CARRYB[21][11] , \CARRYB[21][10] , \CARRYB[21][9] ,
         \CARRYB[21][8] , \CARRYB[21][7] , \CARRYB[21][6] , \CARRYB[21][5] ,
         \CARRYB[21][4] , \CARRYB[21][3] , \CARRYB[21][2] , \CARRYB[21][1] ,
         \CARRYB[21][0] , \CARRYB[20][22] , \CARRYB[20][21] , \CARRYB[20][20] ,
         \CARRYB[20][19] , \CARRYB[20][18] , \CARRYB[20][17] ,
         \CARRYB[20][16] , \CARRYB[20][15] , \CARRYB[20][14] ,
         \CARRYB[20][13] , \CARRYB[20][12] , \CARRYB[20][11] ,
         \CARRYB[20][10] , \CARRYB[20][9] , \CARRYB[20][8] , \CARRYB[20][7] ,
         \CARRYB[20][6] , \CARRYB[20][5] , \CARRYB[20][4] , \CARRYB[20][3] ,
         \CARRYB[20][2] , \CARRYB[20][1] , \CARRYB[20][0] , \CARRYB[19][22] ,
         \CARRYB[19][21] , \CARRYB[19][20] , \CARRYB[19][19] ,
         \CARRYB[19][18] , \CARRYB[19][17] , \CARRYB[19][16] ,
         \CARRYB[19][15] , \CARRYB[19][14] , \CARRYB[19][13] ,
         \CARRYB[19][12] , \CARRYB[19][11] , \CARRYB[19][10] , \CARRYB[19][9] ,
         \CARRYB[19][8] , \CARRYB[19][7] , \CARRYB[19][6] , \CARRYB[19][5] ,
         \CARRYB[19][4] , \CARRYB[19][3] , \CARRYB[19][2] , \CARRYB[19][1] ,
         \CARRYB[19][0] , \CARRYB[18][22] , \CARRYB[18][21] , \CARRYB[18][20] ,
         \CARRYB[18][19] , \CARRYB[18][18] , \CARRYB[18][17] ,
         \CARRYB[18][16] , \CARRYB[18][15] , \CARRYB[18][14] ,
         \CARRYB[18][13] , \CARRYB[18][12] , \CARRYB[18][11] ,
         \CARRYB[18][10] , \CARRYB[18][9] , \CARRYB[18][8] , \CARRYB[18][7] ,
         \CARRYB[18][6] , \CARRYB[18][5] , \CARRYB[18][4] , \CARRYB[18][3] ,
         \CARRYB[18][2] , \CARRYB[18][1] , \CARRYB[18][0] , \CARRYB[17][22] ,
         \CARRYB[17][21] , \CARRYB[17][20] , \CARRYB[17][19] ,
         \CARRYB[17][18] , \CARRYB[17][17] , \CARRYB[17][16] ,
         \CARRYB[17][15] , \CARRYB[17][14] , \CARRYB[17][13] ,
         \CARRYB[17][12] , \CARRYB[17][11] , \CARRYB[17][10] , \CARRYB[17][9] ,
         \CARRYB[17][8] , \CARRYB[17][7] , \CARRYB[17][6] , \CARRYB[17][5] ,
         \CARRYB[17][4] , \CARRYB[17][3] , \CARRYB[17][2] , \CARRYB[17][1] ,
         \CARRYB[17][0] , \CARRYB[16][22] , \CARRYB[16][21] , \CARRYB[16][20] ,
         \CARRYB[16][19] , \CARRYB[16][18] , \CARRYB[16][17] ,
         \CARRYB[16][16] , \CARRYB[16][15] , \CARRYB[16][14] ,
         \CARRYB[16][13] , \CARRYB[16][12] , \CARRYB[16][11] ,
         \CARRYB[16][10] , \CARRYB[16][9] , \CARRYB[16][8] , \CARRYB[16][7] ,
         \CARRYB[16][6] , \CARRYB[16][5] , \CARRYB[16][4] , \CARRYB[16][3] ,
         \CARRYB[16][2] , \CARRYB[16][1] , \CARRYB[16][0] , \CARRYB[15][22] ,
         \CARRYB[15][21] , \CARRYB[15][20] , \CARRYB[15][19] ,
         \CARRYB[15][18] , \CARRYB[15][17] , \CARRYB[15][16] ,
         \CARRYB[15][15] , \CARRYB[15][14] , \CARRYB[15][13] ,
         \CARRYB[15][12] , \CARRYB[15][11] , \CARRYB[15][10] , \CARRYB[15][9] ,
         \CARRYB[15][8] , \CARRYB[15][7] , \CARRYB[15][6] , \CARRYB[15][5] ,
         \CARRYB[15][4] , \CARRYB[15][3] , \CARRYB[15][2] , \CARRYB[15][1] ,
         \CARRYB[15][0] , \CARRYB[14][22] , \CARRYB[14][21] , \CARRYB[14][20] ,
         \CARRYB[14][19] , \CARRYB[14][18] , \CARRYB[14][17] ,
         \CARRYB[14][16] , \CARRYB[14][15] , \CARRYB[14][14] ,
         \CARRYB[14][13] , \CARRYB[14][12] , \CARRYB[14][11] ,
         \CARRYB[14][10] , \CARRYB[14][9] , \CARRYB[14][8] , \CARRYB[14][7] ,
         \CARRYB[14][6] , \CARRYB[14][5] , \CARRYB[14][4] , \CARRYB[14][3] ,
         \CARRYB[14][2] , \CARRYB[14][1] , \CARRYB[14][0] , \CARRYB[13][22] ,
         \CARRYB[13][21] , \CARRYB[13][20] , \CARRYB[13][19] ,
         \CARRYB[13][18] , \CARRYB[13][17] , \CARRYB[13][16] ,
         \CARRYB[13][15] , \CARRYB[13][14] , \CARRYB[13][13] ,
         \CARRYB[13][12] , \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] ,
         \CARRYB[13][8] , \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] ,
         \CARRYB[13][4] , \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] ,
         \CARRYB[13][0] , \CARRYB[12][22] , \CARRYB[12][21] , \CARRYB[12][20] ,
         \CARRYB[12][19] , \CARRYB[12][18] , \CARRYB[12][17] ,
         \CARRYB[12][16] , \CARRYB[12][15] , \CARRYB[12][14] ,
         \CARRYB[12][13] , \CARRYB[12][12] , \CARRYB[12][11] ,
         \CARRYB[12][10] , \CARRYB[12][9] , \CARRYB[12][8] , \CARRYB[12][7] ,
         \CARRYB[12][6] , \CARRYB[12][5] , \CARRYB[12][4] , \CARRYB[12][3] ,
         \CARRYB[12][2] , \CARRYB[12][1] , \CARRYB[12][0] , \CARRYB[11][22] ,
         \CARRYB[11][21] , \CARRYB[11][20] , \CARRYB[11][19] ,
         \CARRYB[11][18] , \CARRYB[11][17] , \CARRYB[11][16] ,
         \CARRYB[11][15] , \CARRYB[11][14] , \CARRYB[11][13] ,
         \CARRYB[11][12] , \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] ,
         \CARRYB[11][8] , \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] ,
         \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] ,
         \CARRYB[11][0] , \CARRYB[10][22] , \CARRYB[10][21] , \CARRYB[10][20] ,
         \CARRYB[10][19] , \CARRYB[10][18] , \CARRYB[10][17] ,
         \CARRYB[10][16] , \CARRYB[10][15] , \CARRYB[10][14] ,
         \CARRYB[10][13] , \CARRYB[10][12] , \CARRYB[10][11] ,
         \CARRYB[10][10] , \CARRYB[10][9] , \CARRYB[10][8] , \CARRYB[10][7] ,
         \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] , \CARRYB[10][3] ,
         \CARRYB[10][2] , \CARRYB[10][1] , \CARRYB[10][0] , \CARRYB[9][22] ,
         \CARRYB[9][21] , \CARRYB[9][20] , \CARRYB[9][19] , \CARRYB[9][18] ,
         \CARRYB[9][17] , \CARRYB[9][16] , \CARRYB[9][15] , \CARRYB[9][14] ,
         \CARRYB[9][13] , \CARRYB[9][12] , \CARRYB[9][11] , \CARRYB[9][10] ,
         \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] ,
         \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] ,
         \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][22] , \CARRYB[8][21] ,
         \CARRYB[8][20] , \CARRYB[8][19] , \CARRYB[8][18] , \CARRYB[8][17] ,
         \CARRYB[8][16] , \CARRYB[8][15] , \CARRYB[8][14] , \CARRYB[8][13] ,
         \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] ,
         \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] ,
         \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] ,
         \CARRYB[8][0] , \CARRYB[7][22] , \CARRYB[7][21] , \CARRYB[7][20] ,
         \CARRYB[7][19] , \CARRYB[7][18] , \CARRYB[7][17] , \CARRYB[7][16] ,
         \CARRYB[7][15] , \CARRYB[7][14] , \CARRYB[7][13] , \CARRYB[7][12] ,
         \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] , \CARRYB[7][8] ,
         \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] , \CARRYB[7][4] ,
         \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] , \CARRYB[7][0] ,
         \CARRYB[6][22] , \CARRYB[6][21] , \CARRYB[6][20] , \CARRYB[6][19] ,
         \CARRYB[6][18] , \CARRYB[6][17] , \CARRYB[6][16] , \CARRYB[6][15] ,
         \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] , \CARRYB[6][11] ,
         \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] , \CARRYB[6][7] ,
         \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] , \CARRYB[6][3] ,
         \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][22] ,
         \CARRYB[5][21] , \CARRYB[5][20] , \CARRYB[5][19] , \CARRYB[5][18] ,
         \CARRYB[5][17] , \CARRYB[5][16] , \CARRYB[5][15] , \CARRYB[5][14] ,
         \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] ,
         \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] ,
         \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] ,
         \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][22] , \CARRYB[4][21] ,
         \CARRYB[4][20] , \CARRYB[4][19] , \CARRYB[4][18] , \CARRYB[4][17] ,
         \CARRYB[4][16] , \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] ,
         \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][22] , \CARRYB[3][21] , \CARRYB[3][20] ,
         \CARRYB[3][19] , \CARRYB[3][18] , \CARRYB[3][17] , \CARRYB[3][16] ,
         \CARRYB[3][15] , \CARRYB[3][14] , \CARRYB[3][13] , \CARRYB[3][12] ,
         \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] , \CARRYB[3][8] ,
         \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] ,
         \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] ,
         \CARRYB[2][22] , \CARRYB[2][21] , \CARRYB[2][20] , \CARRYB[2][19] ,
         \CARRYB[2][18] , \CARRYB[2][17] , \CARRYB[2][16] , \CARRYB[2][15] ,
         \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] , \CARRYB[2][11] ,
         \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] ,
         \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] ,
         \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] , \CARRYB[1][22] ,
         \CARRYB[1][21] , \CARRYB[1][20] , \CARRYB[1][19] , \CARRYB[1][18] ,
         \CARRYB[1][17] , \CARRYB[1][16] , \CARRYB[1][15] , \CARRYB[1][14] ,
         \CARRYB[1][13] , \CARRYB[1][12] , \CARRYB[1][11] , \CARRYB[1][10] ,
         \CARRYB[1][9] , \CARRYB[1][8] , \CARRYB[1][7] , \CARRYB[1][6] ,
         \CARRYB[1][5] , \CARRYB[1][4] , \CARRYB[1][3] , \CARRYB[1][2] ,
         \CARRYB[1][1] , \CARRYB[1][0] , \SUMB[23][22] , \SUMB[23][21] ,
         \SUMB[23][20] , \SUMB[23][19] , \SUMB[23][18] , \SUMB[23][17] ,
         \SUMB[23][16] , \SUMB[23][15] , \SUMB[23][14] , \SUMB[23][13] ,
         \SUMB[23][12] , \SUMB[23][11] , \SUMB[23][10] , \SUMB[23][9] ,
         \SUMB[23][8] , \SUMB[23][7] , \SUMB[23][6] , \SUMB[23][5] ,
         \SUMB[23][4] , \SUMB[23][3] , \SUMB[23][2] , \SUMB[23][1] ,
         \SUMB[23][0] , \SUMB[22][22] , \SUMB[22][21] , \SUMB[22][20] ,
         \SUMB[22][19] , \SUMB[22][18] , \SUMB[22][17] , \SUMB[22][16] ,
         \SUMB[22][15] , \SUMB[22][14] , \SUMB[22][13] , \SUMB[22][12] ,
         \SUMB[22][11] , \SUMB[22][10] , \SUMB[22][9] , \SUMB[22][8] ,
         \SUMB[22][7] , \SUMB[22][6] , \SUMB[22][5] , \SUMB[22][4] ,
         \SUMB[22][3] , \SUMB[22][2] , \SUMB[22][1] , \SUMB[21][22] ,
         \SUMB[21][21] , \SUMB[21][20] , \SUMB[21][19] , \SUMB[21][18] ,
         \SUMB[21][17] , \SUMB[21][16] , \SUMB[21][15] , \SUMB[21][14] ,
         \SUMB[21][13] , \SUMB[21][12] , \SUMB[21][11] , \SUMB[21][10] ,
         \SUMB[21][9] , \SUMB[21][8] , \SUMB[21][7] , \SUMB[21][6] ,
         \SUMB[21][5] , \SUMB[21][4] , \SUMB[21][3] , \SUMB[21][2] ,
         \SUMB[21][1] , \SUMB[20][22] , \SUMB[20][21] , \SUMB[20][20] ,
         \SUMB[20][19] , \SUMB[20][18] , \SUMB[20][17] , \SUMB[20][16] ,
         \SUMB[20][15] , \SUMB[20][14] , \SUMB[20][13] , \SUMB[20][12] ,
         \SUMB[20][11] , \SUMB[20][10] , \SUMB[20][9] , \SUMB[20][8] ,
         \SUMB[20][7] , \SUMB[20][6] , \SUMB[20][5] , \SUMB[20][4] ,
         \SUMB[20][3] , \SUMB[20][2] , \SUMB[20][1] , \SUMB[19][22] ,
         \SUMB[19][21] , \SUMB[19][20] , \SUMB[19][19] , \SUMB[19][18] ,
         \SUMB[19][17] , \SUMB[19][16] , \SUMB[19][15] , \SUMB[19][14] ,
         \SUMB[19][13] , \SUMB[19][12] , \SUMB[19][11] , \SUMB[19][10] ,
         \SUMB[19][9] , \SUMB[19][8] , \SUMB[19][7] , \SUMB[19][6] ,
         \SUMB[19][5] , \SUMB[19][4] , \SUMB[19][3] , \SUMB[19][2] ,
         \SUMB[19][1] , \SUMB[18][22] , \SUMB[18][21] , \SUMB[18][20] ,
         \SUMB[18][19] , \SUMB[18][18] , \SUMB[18][17] , \SUMB[18][16] ,
         \SUMB[18][15] , \SUMB[18][14] , \SUMB[18][13] , \SUMB[18][12] ,
         \SUMB[18][11] , \SUMB[18][10] , \SUMB[18][9] , \SUMB[18][8] ,
         \SUMB[18][7] , \SUMB[18][6] , \SUMB[18][5] , \SUMB[18][4] ,
         \SUMB[18][3] , \SUMB[18][2] , \SUMB[18][1] , \SUMB[17][22] ,
         \SUMB[17][21] , \SUMB[17][20] , \SUMB[17][19] , \SUMB[17][18] ,
         \SUMB[17][17] , \SUMB[17][16] , \SUMB[17][15] , \SUMB[17][14] ,
         \SUMB[17][13] , \SUMB[17][12] , \SUMB[17][11] , \SUMB[17][10] ,
         \SUMB[17][9] , \SUMB[17][8] , \SUMB[17][7] , \SUMB[17][6] ,
         \SUMB[17][5] , \SUMB[17][4] , \SUMB[17][3] , \SUMB[17][2] ,
         \SUMB[17][1] , \SUMB[16][22] , \SUMB[16][21] , \SUMB[16][20] ,
         \SUMB[16][19] , \SUMB[16][18] , \SUMB[16][17] , \SUMB[16][16] ,
         \SUMB[16][15] , \SUMB[16][14] , \SUMB[16][13] , \SUMB[16][12] ,
         \SUMB[16][11] , \SUMB[16][10] , \SUMB[16][9] , \SUMB[16][8] ,
         \SUMB[16][7] , \SUMB[16][6] , \SUMB[16][5] , \SUMB[16][4] ,
         \SUMB[16][3] , \SUMB[16][2] , \SUMB[16][1] , \SUMB[15][22] ,
         \SUMB[15][21] , \SUMB[15][20] , \SUMB[15][19] , \SUMB[15][18] ,
         \SUMB[15][17] , \SUMB[15][16] , \SUMB[15][15] , \SUMB[15][14] ,
         \SUMB[15][13] , \SUMB[15][12] , \SUMB[15][11] , \SUMB[15][10] ,
         \SUMB[15][9] , \SUMB[15][8] , \SUMB[15][7] , \SUMB[15][6] ,
         \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] , \SUMB[15][2] ,
         \SUMB[15][1] , \SUMB[14][22] , \SUMB[14][21] , \SUMB[14][20] ,
         \SUMB[14][19] , \SUMB[14][18] , \SUMB[14][17] , \SUMB[14][16] ,
         \SUMB[14][15] , \SUMB[14][14] , \SUMB[14][13] , \SUMB[14][12] ,
         \SUMB[14][11] , \SUMB[14][10] , \SUMB[14][9] , \SUMB[14][8] ,
         \SUMB[14][7] , \SUMB[14][6] , \SUMB[14][5] , \SUMB[14][4] ,
         \SUMB[14][3] , \SUMB[14][2] , \SUMB[14][1] , \SUMB[13][22] ,
         \SUMB[13][21] , \SUMB[13][20] , \SUMB[13][19] , \SUMB[13][18] ,
         \SUMB[13][17] , \SUMB[13][16] , \SUMB[13][15] , \SUMB[13][14] ,
         \SUMB[13][13] , \SUMB[13][12] , \SUMB[13][11] , \SUMB[13][10] ,
         \SUMB[13][9] , \SUMB[13][8] , \SUMB[13][7] , \SUMB[13][6] ,
         \SUMB[13][5] , \SUMB[13][4] , \SUMB[13][3] , \SUMB[13][2] ,
         \SUMB[13][1] , \SUMB[12][22] , \SUMB[12][21] , \SUMB[12][20] ,
         \SUMB[12][19] , \SUMB[12][18] , \SUMB[12][17] , \SUMB[12][16] ,
         \SUMB[12][15] , \SUMB[12][14] , \SUMB[12][13] , \SUMB[12][12] ,
         \SUMB[12][11] , \SUMB[12][10] , \SUMB[12][9] , \SUMB[12][8] ,
         \SUMB[12][7] , \SUMB[12][6] , \SUMB[12][5] , \SUMB[12][4] ,
         \SUMB[12][3] , \SUMB[12][2] , \SUMB[12][1] , \SUMB[11][22] ,
         \SUMB[11][21] , \SUMB[11][20] , \SUMB[11][19] , \SUMB[11][18] ,
         \SUMB[11][17] , \SUMB[11][16] , \SUMB[11][15] , \SUMB[11][14] ,
         \SUMB[11][13] , \SUMB[11][12] , \SUMB[11][11] , \SUMB[11][10] ,
         \SUMB[11][9] , \SUMB[11][8] , \SUMB[11][7] , \SUMB[11][6] ,
         \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][3] , \SUMB[11][2] ,
         \SUMB[11][1] , \SUMB[10][22] , \SUMB[10][21] , \SUMB[10][20] ,
         \SUMB[10][19] , \SUMB[10][18] , \SUMB[10][17] , \SUMB[10][16] ,
         \SUMB[10][15] , \SUMB[10][14] , \SUMB[10][13] , \SUMB[10][12] ,
         \SUMB[10][11] , \SUMB[10][10] , \SUMB[10][9] , \SUMB[10][8] ,
         \SUMB[10][7] , \SUMB[10][6] , \SUMB[10][5] , \SUMB[10][4] ,
         \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] , \SUMB[9][22] ,
         \SUMB[9][21] , \SUMB[9][20] , \SUMB[9][19] , \SUMB[9][18] ,
         \SUMB[9][17] , \SUMB[9][16] , \SUMB[9][15] , \SUMB[9][14] ,
         \SUMB[9][13] , \SUMB[9][12] , \SUMB[9][11] , \SUMB[9][10] ,
         \SUMB[9][9] , \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] ,
         \SUMB[9][4] , \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][22] ,
         \SUMB[8][21] , \SUMB[8][20] , \SUMB[8][19] , \SUMB[8][18] ,
         \SUMB[8][17] , \SUMB[8][16] , \SUMB[8][15] , \SUMB[8][14] ,
         \SUMB[8][13] , \SUMB[8][12] , \SUMB[8][11] , \SUMB[8][10] ,
         \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] ,
         \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][22] ,
         \SUMB[7][21] , \SUMB[7][20] , \SUMB[7][19] , \SUMB[7][18] ,
         \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] , \SUMB[7][14] ,
         \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] ,
         \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] ,
         \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][22] ,
         \SUMB[6][21] , \SUMB[6][20] , \SUMB[6][19] , \SUMB[6][18] ,
         \SUMB[6][17] , \SUMB[6][16] , \SUMB[6][15] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][22] ,
         \SUMB[5][21] , \SUMB[5][20] , \SUMB[5][19] , \SUMB[5][18] ,
         \SUMB[5][17] , \SUMB[5][16] , \SUMB[5][15] , \SUMB[5][14] ,
         \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] ,
         \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][22] ,
         \SUMB[4][21] , \SUMB[4][20] , \SUMB[4][19] , \SUMB[4][18] ,
         \SUMB[4][17] , \SUMB[4][16] , \SUMB[4][15] , \SUMB[4][14] ,
         \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][22] ,
         \SUMB[3][21] , \SUMB[3][20] , \SUMB[3][19] , \SUMB[3][18] ,
         \SUMB[3][17] , \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][22] ,
         \SUMB[2][21] , \SUMB[2][20] , \SUMB[2][19] , \SUMB[2][18] ,
         \SUMB[2][17] , \SUMB[2][16] , \SUMB[2][15] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][22] ,
         \SUMB[1][21] , \SUMB[1][20] , \SUMB[1][19] , \SUMB[1][18] ,
         \SUMB[1][17] , \SUMB[1][16] , \SUMB[1][15] , \SUMB[1][14] ,
         \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] , \SUMB[1][10] ,
         \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] ,
         \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , \A1[43] ,
         \A1[42] , \A1[41] , \A1[40] , \A1[39] , \A1[38] , \A1[37] , \A1[36] ,
         \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] ,
         \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] ,
         \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] ,
         \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] ,
         \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] ,
         \A2[44] , \A2[43] , \A2[42] , \A2[41] , \A2[40] , \A2[39] , \A2[38] ,
         \A2[37] , \A2[36] , \A2[35] , \A2[34] , \A2[33] , \A2[32] , \A2[31] ,
         \A2[30] , \A2[29] , \A2[28] , \A2[27] , \A2[26] , \A2[25] , \A2[24] ,
         \A2[23] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95;
  assign \ab[23][22]  = B[22];
  assign \ab[23][21]  = B[21];
  assign \ab[23][20]  = B[20];
  assign \ab[23][19]  = B[19];
  assign \ab[23][18]  = B[18];
  assign \ab[23][17]  = B[17];
  assign \ab[23][16]  = B[16];
  assign \ab[23][15]  = B[15];
  assign \ab[23][14]  = B[14];
  assign \ab[23][13]  = B[13];
  assign \ab[23][12]  = B[12];
  assign \ab[23][11]  = B[11];
  assign \ab[23][10]  = B[10];
  assign \ab[23][9]  = B[9];
  assign \ab[23][8]  = B[8];
  assign \ab[23][7]  = B[7];
  assign \ab[23][6]  = B[6];
  assign \ab[23][5]  = B[5];
  assign \ab[23][4]  = B[4];
  assign \ab[23][3]  = B[3];
  assign \ab[23][2]  = B[2];
  assign \ab[23][1]  = B[1];
  assign \ab[23][0]  = B[0];
  assign \ab[22][23]  = A[22];
  assign \ab[21][23]  = A[21];
  assign \ab[20][23]  = A[20];
  assign \ab[19][23]  = A[19];
  assign \ab[18][23]  = A[18];
  assign \ab[17][23]  = A[17];
  assign \ab[16][23]  = A[16];
  assign \ab[15][23]  = A[15];
  assign \ab[14][23]  = A[14];
  assign \ab[13][23]  = A[13];
  assign \ab[12][23]  = A[12];
  assign \ab[11][23]  = A[11];
  assign \ab[10][23]  = A[10];
  assign \ab[9][23]  = A[9];
  assign \ab[8][23]  = A[8];
  assign \ab[7][23]  = A[7];
  assign \ab[6][23]  = A[6];
  assign \ab[5][23]  = A[5];
  assign \ab[4][23]  = A[4];
  assign \ab[3][23]  = A[3];
  assign \ab[2][23]  = A[2];
  assign \ab[1][23]  = A[1];
  assign \ab[0][23]  = A[0];

  FPU_CAL_DW01_add_2 FS_1 ( .A({1'b0, n95, \A1[43] , \A1[42] , \A1[41] , 
        \A1[40] , \A1[39] , \A1[38] , \A1[37] , \A1[36] , \A1[35] , \A1[34] , 
        \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] , \A1[27] , 
        \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \SUMB[23][0] , 
        \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , 
        \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , 
        \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({
        \CARRYB[23][22] , \A2[44] , \A2[43] , \A2[42] , \A2[41] , \A2[40] , 
        \A2[39] , \A2[38] , \A2[37] , \A2[36] , \A2[35] , \A2[34] , \A2[33] , 
        \A2[32] , \A2[31] , \A2[30] , \A2[29] , \A2[28] , \A2[27] , \A2[26] , 
        \A2[25] , \A2[24] , \A2[23] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM(PRODUCT[47:2]) );
  FADDX1_RVT S2_22_20 ( .A(\ab[22][20] ), .B(\CARRYB[21][20] ), .CI(
        \SUMB[21][21] ), .CO(\CARRYB[22][20] ), .S(\SUMB[22][20] ) );
  FADDX1_RVT S2_21_20 ( .A(\ab[21][20] ), .B(\CARRYB[20][20] ), .CI(
        \SUMB[20][21] ), .CO(\CARRYB[21][20] ), .S(\SUMB[21][20] ) );
  FADDX1_RVT S2_20_20 ( .A(\ab[20][20] ), .B(\CARRYB[19][20] ), .CI(
        \SUMB[19][21] ), .CO(\CARRYB[20][20] ), .S(\SUMB[20][20] ) );
  FADDX1_RVT S2_22_18 ( .A(\ab[22][18] ), .B(\CARRYB[21][18] ), .CI(
        \SUMB[21][19] ), .CO(\CARRYB[22][18] ), .S(\SUMB[22][18] ) );
  FADDX1_RVT S2_22_19 ( .A(\ab[22][19] ), .B(\CARRYB[21][19] ), .CI(
        \SUMB[21][20] ), .CO(\CARRYB[22][19] ), .S(\SUMB[22][19] ) );
  FADDX1_RVT S2_21_19 ( .A(\ab[21][19] ), .B(\CARRYB[20][19] ), .CI(
        \SUMB[20][20] ), .CO(\CARRYB[21][19] ), .S(\SUMB[21][19] ) );
  FADDX1_RVT S3_22_22 ( .A(\ab[22][22] ), .B(\CARRYB[21][22] ), .CI(n91), .CO(
        \CARRYB[22][22] ), .S(\SUMB[22][22] ) );
  FADDX1_RVT S2_19_21 ( .A(\ab[19][21] ), .B(\CARRYB[18][21] ), .CI(
        \SUMB[18][22] ), .CO(\CARRYB[19][21] ), .S(\SUMB[19][21] ) );
  FADDX1_RVT S2_22_21 ( .A(\ab[22][21] ), .B(\CARRYB[21][21] ), .CI(
        \SUMB[21][22] ), .CO(\CARRYB[22][21] ), .S(\SUMB[22][21] ) );
  FADDX1_RVT S2_20_21 ( .A(\ab[20][21] ), .B(\CARRYB[19][21] ), .CI(
        \SUMB[19][22] ), .CO(\CARRYB[20][21] ), .S(\SUMB[20][21] ) );
  FADDX1_RVT S2_21_21 ( .A(\ab[21][21] ), .B(\CARRYB[20][21] ), .CI(
        \SUMB[20][22] ), .CO(\CARRYB[21][21] ), .S(\SUMB[21][21] ) );
  FADDX1_RVT S4_20 ( .A(n43), .B(\CARRYB[22][20] ), .CI(\SUMB[22][21] ), .CO(
        \CARRYB[23][20] ), .S(\SUMB[23][20] ) );
  FADDX1_RVT S4_17 ( .A(n37), .B(\CARRYB[22][17] ), .CI(\SUMB[22][18] ), .CO(
        \CARRYB[23][17] ), .S(\SUMB[23][17] ) );
  FADDX1_RVT S5_22 ( .A(n47), .B(\CARRYB[22][22] ), .CI(n93), .CO(
        \CARRYB[23][22] ), .S(\SUMB[23][22] ) );
  FADDX1_RVT S4_18 ( .A(n39), .B(\CARRYB[22][18] ), .CI(\SUMB[22][19] ), .CO(
        \CARRYB[23][18] ), .S(\SUMB[23][18] ) );
  FADDX1_RVT S4_21 ( .A(n45), .B(\CARRYB[22][21] ), .CI(\SUMB[22][22] ), .CO(
        \CARRYB[23][21] ), .S(\SUMB[23][21] ) );
  FADDX1_RVT S4_19 ( .A(n41), .B(\CARRYB[22][19] ), .CI(\SUMB[22][20] ), .CO(
        \CARRYB[23][19] ), .S(\SUMB[23][19] ) );
  FADDX1_RVT S3_18_22 ( .A(\ab[18][22] ), .B(\CARRYB[17][22] ), .CI(n83), .CO(
        \CARRYB[18][22] ), .S(\SUMB[18][22] ) );
  FADDX1_RVT S3_21_22 ( .A(\ab[21][22] ), .B(\CARRYB[20][22] ), .CI(n89), .CO(
        \CARRYB[21][22] ), .S(\SUMB[21][22] ) );
  FADDX1_RVT S3_19_22 ( .A(\ab[19][22] ), .B(\CARRYB[18][22] ), .CI(n85), .CO(
        \CARRYB[19][22] ), .S(\SUMB[19][22] ) );
  FADDX1_RVT S3_20_22 ( .A(\ab[20][22] ), .B(\CARRYB[19][22] ), .CI(n87), .CO(
        \CARRYB[20][22] ), .S(\SUMB[20][22] ) );
  FADDX1_RVT S2_22_1 ( .A(\ab[22][1] ), .B(\CARRYB[21][1] ), .CI(\SUMB[21][2] ), .CO(\CARRYB[22][1] ), .S(\SUMB[22][1] ) );
  FADDX1_RVT S2_21_1 ( .A(\ab[21][1] ), .B(\CARRYB[20][1] ), .CI(\SUMB[20][2] ), .CO(\CARRYB[21][1] ), .S(\SUMB[21][1] ) );
  FADDX1_RVT S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), 
        .CO(\CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FADDX1_RVT S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), 
        .CO(\CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FADDX1_RVT S1_22_0 ( .A(\ab[22][0] ), .B(\CARRYB[21][0] ), .CI(\SUMB[21][1] ), .CO(\CARRYB[22][0] ), .S(\A1[20] ) );
  FADDX1_RVT S1_21_0 ( .A(\ab[21][0] ), .B(\CARRYB[20][0] ), .CI(\SUMB[20][1] ), .CO(\CARRYB[21][0] ), .S(\A1[19] ) );
  FADDX1_RVT S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), 
        .CO(\CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FADDX1_RVT S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), 
        .CO(\CARRYB[10][0] ), .S(\A1[8] ) );
  FADDX1_RVT S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), 
        .CO(\CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FADDX1_RVT S2_16_1 ( .A(\ab[16][1] ), .B(\CARRYB[15][1] ), .CI(\SUMB[15][2] ), .CO(\CARRYB[16][1] ), .S(\SUMB[16][1] ) );
  FADDX1_RVT S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FADDX1_RVT S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), 
        .CO(\CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FADDX1_RVT S2_17_1 ( .A(\ab[17][1] ), .B(\CARRYB[16][1] ), .CI(\SUMB[16][2] ), .CO(\CARRYB[17][1] ), .S(\SUMB[17][1] ) );
  FADDX1_RVT S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), 
        .CO(\CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FADDX1_RVT S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FADDX1_RVT S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FADDX1_RVT S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), 
        .CO(\CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FADDX1_RVT S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), 
        .CO(\CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FADDX1_RVT S2_20_1 ( .A(\ab[20][1] ), .B(\CARRYB[19][1] ), .CI(\SUMB[19][2] ), .CO(\CARRYB[20][1] ), .S(\SUMB[20][1] ) );
  FADDX1_RVT S2_18_1 ( .A(\ab[18][1] ), .B(\CARRYB[17][1] ), .CI(\SUMB[17][2] ), .CO(\CARRYB[18][1] ), .S(\SUMB[18][1] ) );
  FADDX1_RVT S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), 
        .CO(\CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FADDX1_RVT S2_15_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), .CO(\CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FADDX1_RVT S2_22_2 ( .A(\ab[22][2] ), .B(\CARRYB[21][2] ), .CI(\SUMB[21][3] ), .CO(\CARRYB[22][2] ), .S(\SUMB[22][2] ) );
  FADDX1_RVT S2_21_2 ( .A(\ab[21][2] ), .B(\CARRYB[20][2] ), .CI(\SUMB[20][3] ), .CO(\CARRYB[21][2] ), .S(\SUMB[21][2] ) );
  FADDX1_RVT S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), 
        .CO(\CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FADDX1_RVT S2_19_1 ( .A(\ab[19][1] ), .B(\CARRYB[18][1] ), .CI(\SUMB[18][2] ), .CO(\CARRYB[19][1] ), .S(\SUMB[19][1] ) );
  FADDX1_RVT S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), 
        .CO(\CARRYB[2][0] ), .S(\A1[0] ) );
  FADDX1_RVT S2_2_18 ( .A(\ab[2][18] ), .B(\CARRYB[1][18] ), .CI(\SUMB[1][19] ), .CO(\CARRYB[2][18] ), .S(\SUMB[2][18] ) );
  FADDX1_RVT S2_22_16 ( .A(\ab[22][16] ), .B(\CARRYB[21][16] ), .CI(
        \SUMB[21][17] ), .CO(\CARRYB[22][16] ), .S(\SUMB[22][16] ) );
  FADDX1_RVT S2_21_16 ( .A(\ab[21][16] ), .B(\CARRYB[20][16] ), .CI(
        \SUMB[20][17] ), .CO(\CARRYB[21][16] ), .S(\SUMB[21][16] ) );
  FADDX1_RVT S2_20_16 ( .A(\ab[20][16] ), .B(\CARRYB[19][16] ), .CI(
        \SUMB[19][17] ), .CO(\CARRYB[20][16] ), .S(\SUMB[20][16] ) );
  FADDX1_RVT S2_19_16 ( .A(\ab[19][16] ), .B(\CARRYB[18][16] ), .CI(
        \SUMB[18][17] ), .CO(\CARRYB[19][16] ), .S(\SUMB[19][16] ) );
  FADDX1_RVT S2_18_16 ( .A(\ab[18][16] ), .B(\CARRYB[17][16] ), .CI(
        \SUMB[17][17] ), .CO(\CARRYB[18][16] ), .S(\SUMB[18][16] ) );
  FADDX1_RVT S2_22_6 ( .A(\ab[22][6] ), .B(\CARRYB[21][6] ), .CI(\SUMB[21][7] ), .CO(\CARRYB[22][6] ), .S(\SUMB[22][6] ) );
  FADDX1_RVT S2_17_16 ( .A(\ab[17][16] ), .B(\CARRYB[16][16] ), .CI(
        \SUMB[16][17] ), .CO(\CARRYB[17][16] ), .S(\SUMB[17][16] ) );
  FADDX1_RVT S2_21_6 ( .A(\ab[21][6] ), .B(\CARRYB[20][6] ), .CI(\SUMB[20][7] ), .CO(\CARRYB[21][6] ), .S(\SUMB[21][6] ) );
  FADDX1_RVT S2_20_6 ( .A(\ab[20][6] ), .B(\CARRYB[19][6] ), .CI(\SUMB[19][7] ), .CO(\CARRYB[20][6] ), .S(\SUMB[20][6] ) );
  FADDX1_RVT S2_16_16 ( .A(\ab[16][16] ), .B(\CARRYB[15][16] ), .CI(
        \SUMB[15][17] ), .CO(\CARRYB[16][16] ), .S(\SUMB[16][16] ) );
  FADDX1_RVT S2_15_16 ( .A(\ab[15][16] ), .B(\CARRYB[14][16] ), .CI(
        \SUMB[14][17] ), .CO(\CARRYB[15][16] ), .S(\SUMB[15][16] ) );
  FADDX1_RVT S2_19_6 ( .A(\ab[19][6] ), .B(\CARRYB[18][6] ), .CI(\SUMB[18][7] ), .CO(\CARRYB[19][6] ), .S(\SUMB[19][6] ) );
  FADDX1_RVT S2_14_16 ( .A(\ab[14][16] ), .B(\CARRYB[13][16] ), .CI(
        \SUMB[13][17] ), .CO(\CARRYB[14][16] ), .S(\SUMB[14][16] ) );
  FADDX1_RVT S2_18_6 ( .A(\ab[18][6] ), .B(\CARRYB[17][6] ), .CI(\SUMB[17][7] ), .CO(\CARRYB[18][6] ), .S(\SUMB[18][6] ) );
  FADDX1_RVT S2_17_6 ( .A(\ab[17][6] ), .B(\CARRYB[16][6] ), .CI(\SUMB[16][7] ), .CO(\CARRYB[17][6] ), .S(\SUMB[17][6] ) );
  FADDX1_RVT S2_13_16 ( .A(\ab[13][16] ), .B(\CARRYB[12][16] ), .CI(
        \SUMB[12][17] ), .CO(\CARRYB[13][16] ), .S(\SUMB[13][16] ) );
  FADDX1_RVT S2_16_6 ( .A(\ab[16][6] ), .B(\CARRYB[15][6] ), .CI(\SUMB[15][7] ), .CO(\CARRYB[16][6] ), .S(\SUMB[16][6] ) );
  FADDX1_RVT S2_12_16 ( .A(\ab[12][16] ), .B(\CARRYB[11][16] ), .CI(
        \SUMB[11][17] ), .CO(\CARRYB[12][16] ), .S(\SUMB[12][16] ) );
  FADDX1_RVT S2_15_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), .CO(\CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FADDX1_RVT S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FADDX1_RVT S2_10_16 ( .A(\ab[10][16] ), .B(\CARRYB[9][16] ), .CI(
        \SUMB[9][17] ), .CO(\CARRYB[10][16] ), .S(\SUMB[10][16] ) );
  FADDX1_RVT S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FADDX1_RVT S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FADDX1_RVT S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), 
        .CO(\CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FADDX1_RVT S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), 
        .CO(\CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FADDX1_RVT S2_8_16 ( .A(\ab[8][16] ), .B(\CARRYB[7][16] ), .CI(\SUMB[7][17] ), .CO(\CARRYB[8][16] ), .S(\SUMB[8][16] ) );
  FADDX1_RVT S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), 
        .CO(\CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FADDX1_RVT S2_7_16 ( .A(\ab[7][16] ), .B(\CARRYB[6][16] ), .CI(\SUMB[6][17] ), .CO(\CARRYB[7][16] ), .S(\SUMB[7][16] ) );
  FADDX1_RVT S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), 
        .CO(\CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FADDX1_RVT S2_6_16 ( .A(\ab[6][16] ), .B(\CARRYB[5][16] ), .CI(\SUMB[5][17] ), .CO(\CARRYB[6][16] ), .S(\SUMB[6][16] ) );
  FADDX1_RVT S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), 
        .CO(\CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FADDX1_RVT S2_5_16 ( .A(\ab[5][16] ), .B(\CARRYB[4][16] ), .CI(\SUMB[4][17] ), .CO(\CARRYB[5][16] ), .S(\SUMB[5][16] ) );
  FADDX1_RVT S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), 
        .CO(\CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FADDX1_RVT S2_4_16 ( .A(\ab[4][16] ), .B(\CARRYB[3][16] ), .CI(\SUMB[3][17] ), .CO(\CARRYB[4][16] ), .S(\SUMB[4][16] ) );
  FADDX1_RVT S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), 
        .CO(\CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FADDX1_RVT S2_3_16 ( .A(\ab[3][16] ), .B(\CARRYB[2][16] ), .CI(\SUMB[2][17] ), .CO(\CARRYB[3][16] ), .S(\SUMB[3][16] ) );
  FADDX1_RVT S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), 
        .CO(\CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FADDX1_RVT S2_2_16 ( .A(\ab[2][16] ), .B(\CARRYB[1][16] ), .CI(\SUMB[1][17] ), .CO(\CARRYB[2][16] ), .S(\SUMB[2][16] ) );
  FADDX1_RVT S2_22_12 ( .A(\ab[22][12] ), .B(\CARRYB[21][12] ), .CI(
        \SUMB[21][13] ), .CO(\CARRYB[22][12] ), .S(\SUMB[22][12] ) );
  FADDX1_RVT S2_21_12 ( .A(\ab[21][12] ), .B(\CARRYB[20][12] ), .CI(
        \SUMB[20][13] ), .CO(\CARRYB[21][12] ), .S(\SUMB[21][12] ) );
  FADDX1_RVT S2_20_12 ( .A(\ab[20][12] ), .B(\CARRYB[19][12] ), .CI(
        \SUMB[19][13] ), .CO(\CARRYB[20][12] ), .S(\SUMB[20][12] ) );
  FADDX1_RVT S2_19_12 ( .A(\ab[19][12] ), .B(\CARRYB[18][12] ), .CI(
        \SUMB[18][13] ), .CO(\CARRYB[19][12] ), .S(\SUMB[19][12] ) );
  FADDX1_RVT S2_18_12 ( .A(\ab[18][12] ), .B(\CARRYB[17][12] ), .CI(
        \SUMB[17][13] ), .CO(\CARRYB[18][12] ), .S(\SUMB[18][12] ) );
  FADDX1_RVT S2_17_12 ( .A(\ab[17][12] ), .B(\CARRYB[16][12] ), .CI(
        \SUMB[16][13] ), .CO(\CARRYB[17][12] ), .S(\SUMB[17][12] ) );
  FADDX1_RVT S2_16_12 ( .A(\ab[16][12] ), .B(\CARRYB[15][12] ), .CI(
        \SUMB[15][13] ), .CO(\CARRYB[16][12] ), .S(\SUMB[16][12] ) );
  FADDX1_RVT S2_15_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(
        \SUMB[14][13] ), .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FADDX1_RVT S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(
        \SUMB[13][13] ), .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FADDX1_RVT S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(
        \SUMB[12][13] ), .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FADDX1_RVT S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(
        \SUMB[11][13] ), .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FADDX1_RVT S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FADDX1_RVT S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FADDX1_RVT S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FADDX1_RVT S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FADDX1_RVT S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FADDX1_RVT S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FADDX1_RVT S2_2_12 ( .A(\ab[2][12] ), .B(\CARRYB[1][12] ), .CI(\SUMB[1][13] ), .CO(\CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FADDX1_RVT S2_19_20 ( .A(\ab[19][20] ), .B(\CARRYB[18][20] ), .CI(
        \SUMB[18][21] ), .CO(\CARRYB[19][20] ), .S(\SUMB[19][20] ) );
  FADDX1_RVT S2_18_20 ( .A(\ab[18][20] ), .B(\CARRYB[17][20] ), .CI(
        \SUMB[17][21] ), .CO(\CARRYB[18][20] ), .S(\SUMB[18][20] ) );
  FADDX1_RVT S2_17_20 ( .A(\ab[17][20] ), .B(\CARRYB[16][20] ), .CI(
        \SUMB[16][21] ), .CO(\CARRYB[17][20] ), .S(\SUMB[17][20] ) );
  FADDX1_RVT S2_16_20 ( .A(\ab[16][20] ), .B(\CARRYB[15][20] ), .CI(
        \SUMB[15][21] ), .CO(\CARRYB[16][20] ), .S(\SUMB[16][20] ) );
  FADDX1_RVT S2_15_20 ( .A(\ab[15][20] ), .B(\CARRYB[14][20] ), .CI(
        \SUMB[14][21] ), .CO(\CARRYB[15][20] ), .S(\SUMB[15][20] ) );
  FADDX1_RVT S2_14_20 ( .A(\ab[14][20] ), .B(\CARRYB[13][20] ), .CI(
        \SUMB[13][21] ), .CO(\CARRYB[14][20] ), .S(\SUMB[14][20] ) );
  FADDX1_RVT S2_13_20 ( .A(\ab[13][20] ), .B(\CARRYB[12][20] ), .CI(
        \SUMB[12][21] ), .CO(\CARRYB[13][20] ), .S(\SUMB[13][20] ) );
  FADDX1_RVT S2_12_20 ( .A(\ab[12][20] ), .B(\CARRYB[11][20] ), .CI(
        \SUMB[11][21] ), .CO(\CARRYB[12][20] ), .S(\SUMB[12][20] ) );
  FADDX1_RVT S2_10_20 ( .A(\ab[10][20] ), .B(\CARRYB[9][20] ), .CI(
        \SUMB[9][21] ), .CO(\CARRYB[10][20] ), .S(\SUMB[10][20] ) );
  FADDX1_RVT S2_8_20 ( .A(\ab[8][20] ), .B(\CARRYB[7][20] ), .CI(\SUMB[7][21] ), .CO(\CARRYB[8][20] ), .S(\SUMB[8][20] ) );
  FADDX1_RVT S2_7_20 ( .A(\ab[7][20] ), .B(\CARRYB[6][20] ), .CI(\SUMB[6][21] ), .CO(\CARRYB[7][20] ), .S(\SUMB[7][20] ) );
  FADDX1_RVT S2_6_20 ( .A(\ab[6][20] ), .B(\CARRYB[5][20] ), .CI(\SUMB[5][21] ), .CO(\CARRYB[6][20] ), .S(\SUMB[6][20] ) );
  FADDX1_RVT S2_5_20 ( .A(\ab[5][20] ), .B(\CARRYB[4][20] ), .CI(\SUMB[4][21] ), .CO(\CARRYB[5][20] ), .S(\SUMB[5][20] ) );
  FADDX1_RVT S2_4_20 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .CI(\SUMB[3][21] ), .CO(\CARRYB[4][20] ), .S(\SUMB[4][20] ) );
  FADDX1_RVT S2_3_20 ( .A(\ab[3][20] ), .B(\CARRYB[2][20] ), .CI(\SUMB[2][21] ), .CO(\CARRYB[3][20] ), .S(\SUMB[3][20] ) );
  FADDX1_RVT S2_2_20 ( .A(\ab[2][20] ), .B(\CARRYB[1][20] ), .CI(\SUMB[1][21] ), .CO(\CARRYB[2][20] ), .S(\SUMB[2][20] ) );
  FADDX1_RVT S2_2_17 ( .A(\ab[2][17] ), .B(\CARRYB[1][17] ), .CI(\SUMB[1][18] ), .CO(\CARRYB[2][17] ), .S(\SUMB[2][17] ) );
  FADDX1_RVT S2_22_4 ( .A(\ab[22][4] ), .B(\CARRYB[21][4] ), .CI(\SUMB[21][5] ), .CO(\CARRYB[22][4] ), .S(\SUMB[22][4] ) );
  FADDX1_RVT S2_22_8 ( .A(\ab[22][8] ), .B(\CARRYB[21][8] ), .CI(\SUMB[21][9] ), .CO(\CARRYB[22][8] ), .S(\SUMB[22][8] ) );
  FADDX1_RVT S2_21_8 ( .A(\ab[21][8] ), .B(\CARRYB[20][8] ), .CI(\SUMB[20][9] ), .CO(\CARRYB[21][8] ), .S(\SUMB[21][8] ) );
  FADDX1_RVT S2_20_8 ( .A(\ab[20][8] ), .B(\CARRYB[19][8] ), .CI(\SUMB[19][9] ), .CO(\CARRYB[20][8] ), .S(\SUMB[20][8] ) );
  FADDX1_RVT S2_19_8 ( .A(\ab[19][8] ), .B(\CARRYB[18][8] ), .CI(\SUMB[18][9] ), .CO(\CARRYB[19][8] ), .S(\SUMB[19][8] ) );
  FADDX1_RVT S2_18_8 ( .A(\ab[18][8] ), .B(\CARRYB[17][8] ), .CI(\SUMB[17][9] ), .CO(\CARRYB[18][8] ), .S(\SUMB[18][8] ) );
  FADDX1_RVT S2_21_4 ( .A(\ab[21][4] ), .B(\CARRYB[20][4] ), .CI(\SUMB[20][5] ), .CO(\CARRYB[21][4] ), .S(\SUMB[21][4] ) );
  FADDX1_RVT S2_20_4 ( .A(\ab[20][4] ), .B(\CARRYB[19][4] ), .CI(\SUMB[19][5] ), .CO(\CARRYB[20][4] ), .S(\SUMB[20][4] ) );
  FADDX1_RVT S2_19_4 ( .A(\ab[19][4] ), .B(\CARRYB[18][4] ), .CI(\SUMB[18][5] ), .CO(\CARRYB[19][4] ), .S(\SUMB[19][4] ) );
  FADDX1_RVT S2_17_8 ( .A(\ab[17][8] ), .B(\CARRYB[16][8] ), .CI(\SUMB[16][9] ), .CO(\CARRYB[17][8] ), .S(\SUMB[17][8] ) );
  FADDX1_RVT S2_16_8 ( .A(\ab[16][8] ), .B(\CARRYB[15][8] ), .CI(\SUMB[15][9] ), .CO(\CARRYB[16][8] ), .S(\SUMB[16][8] ) );
  FADDX1_RVT S2_15_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), .CO(\CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FADDX1_RVT S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FADDX1_RVT S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FADDX1_RVT S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), 
        .CO(\CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FADDX1_RVT S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), 
        .CO(\CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FADDX1_RVT S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), 
        .CO(\CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FADDX1_RVT S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), 
        .CO(\CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FADDX1_RVT S2_22_17 ( .A(\ab[22][17] ), .B(\CARRYB[21][17] ), .CI(
        \SUMB[21][18] ), .CO(\CARRYB[22][17] ), .S(\SUMB[22][17] ) );
  FADDX1_RVT S2_21_17 ( .A(\ab[21][17] ), .B(\CARRYB[20][17] ), .CI(
        \SUMB[20][18] ), .CO(\CARRYB[21][17] ), .S(\SUMB[21][17] ) );
  FADDX1_RVT S2_20_17 ( .A(\ab[20][17] ), .B(\CARRYB[19][17] ), .CI(
        \SUMB[19][18] ), .CO(\CARRYB[20][17] ), .S(\SUMB[20][17] ) );
  FADDX1_RVT S2_19_17 ( .A(\ab[19][17] ), .B(\CARRYB[18][17] ), .CI(
        \SUMB[18][18] ), .CO(\CARRYB[19][17] ), .S(\SUMB[19][17] ) );
  FADDX1_RVT S2_18_17 ( .A(\ab[18][17] ), .B(\CARRYB[17][17] ), .CI(
        \SUMB[17][18] ), .CO(\CARRYB[18][17] ), .S(\SUMB[18][17] ) );
  FADDX1_RVT S2_17_17 ( .A(\ab[17][17] ), .B(\CARRYB[16][17] ), .CI(
        \SUMB[16][18] ), .CO(\CARRYB[17][17] ), .S(\SUMB[17][17] ) );
  FADDX1_RVT S2_22_7 ( .A(\ab[22][7] ), .B(\CARRYB[21][7] ), .CI(\SUMB[21][8] ), .CO(\CARRYB[22][7] ), .S(\SUMB[22][7] ) );
  FADDX1_RVT S2_21_7 ( .A(\ab[21][7] ), .B(\CARRYB[20][7] ), .CI(\SUMB[20][8] ), .CO(\CARRYB[21][7] ), .S(\SUMB[21][7] ) );
  FADDX1_RVT S2_16_17 ( .A(\ab[16][17] ), .B(\CARRYB[15][17] ), .CI(
        \SUMB[15][18] ), .CO(\CARRYB[16][17] ), .S(\SUMB[16][17] ) );
  FADDX1_RVT S2_20_7 ( .A(\ab[20][7] ), .B(\CARRYB[19][7] ), .CI(\SUMB[19][8] ), .CO(\CARRYB[20][7] ), .S(\SUMB[20][7] ) );
  FADDX1_RVT S2_19_7 ( .A(\ab[19][7] ), .B(\CARRYB[18][7] ), .CI(\SUMB[18][8] ), .CO(\CARRYB[19][7] ), .S(\SUMB[19][7] ) );
  FADDX1_RVT S2_22_3 ( .A(\ab[22][3] ), .B(\CARRYB[21][3] ), .CI(\SUMB[21][4] ), .CO(\CARRYB[22][3] ), .S(\SUMB[22][3] ) );
  FADDX1_RVT S2_15_17 ( .A(\ab[15][17] ), .B(\CARRYB[14][17] ), .CI(
        \SUMB[14][18] ), .CO(\CARRYB[15][17] ), .S(\SUMB[15][17] ) );
  FADDX1_RVT S2_21_3 ( .A(\ab[21][3] ), .B(\CARRYB[20][3] ), .CI(\SUMB[20][4] ), .CO(\CARRYB[21][3] ), .S(\SUMB[21][3] ) );
  FADDX1_RVT S2_20_3 ( .A(\ab[20][3] ), .B(\CARRYB[19][3] ), .CI(\SUMB[19][4] ), .CO(\CARRYB[20][3] ), .S(\SUMB[20][3] ) );
  FADDX1_RVT S2_14_17 ( .A(\ab[14][17] ), .B(\CARRYB[13][17] ), .CI(
        \SUMB[13][18] ), .CO(\CARRYB[14][17] ), .S(\SUMB[14][17] ) );
  FADDX1_RVT S2_19_3 ( .A(\ab[19][3] ), .B(\CARRYB[18][3] ), .CI(\SUMB[18][4] ), .CO(\CARRYB[19][3] ), .S(\SUMB[19][3] ) );
  FADDX1_RVT S2_18_3 ( .A(\ab[18][3] ), .B(\CARRYB[17][3] ), .CI(\SUMB[17][4] ), .CO(\CARRYB[18][3] ), .S(\SUMB[18][3] ) );
  FADDX1_RVT S2_18_7 ( .A(\ab[18][7] ), .B(\CARRYB[17][7] ), .CI(\SUMB[17][8] ), .CO(\CARRYB[18][7] ), .S(\SUMB[18][7] ) );
  FADDX1_RVT S2_13_17 ( .A(\ab[13][17] ), .B(\CARRYB[12][17] ), .CI(
        \SUMB[12][18] ), .CO(\CARRYB[13][17] ), .S(\SUMB[13][17] ) );
  FADDX1_RVT S2_17_3 ( .A(\ab[17][3] ), .B(\CARRYB[16][3] ), .CI(\SUMB[16][4] ), .CO(\CARRYB[17][3] ), .S(\SUMB[17][3] ) );
  FADDX1_RVT S2_17_7 ( .A(\ab[17][7] ), .B(\CARRYB[16][7] ), .CI(\SUMB[16][8] ), .CO(\CARRYB[17][7] ), .S(\SUMB[17][7] ) );
  FADDX1_RVT S2_16_3 ( .A(\ab[16][3] ), .B(\CARRYB[15][3] ), .CI(\SUMB[15][4] ), .CO(\CARRYB[16][3] ), .S(\SUMB[16][3] ) );
  FADDX1_RVT S2_16_7 ( .A(\ab[16][7] ), .B(\CARRYB[15][7] ), .CI(\SUMB[15][8] ), .CO(\CARRYB[16][7] ), .S(\SUMB[16][7] ) );
  FADDX1_RVT S2_12_17 ( .A(\ab[12][17] ), .B(\CARRYB[11][17] ), .CI(
        \SUMB[11][18] ), .CO(\CARRYB[12][17] ), .S(\SUMB[12][17] ) );
  FADDX1_RVT S2_15_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), .CO(\CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FADDX1_RVT S2_15_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), .CO(\CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FADDX1_RVT S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FADDX1_RVT S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FADDX1_RVT S2_10_17 ( .A(\ab[10][17] ), .B(\CARRYB[9][17] ), .CI(
        \SUMB[9][18] ), .CO(\CARRYB[10][17] ), .S(\SUMB[10][17] ) );
  FADDX1_RVT S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FADDX1_RVT S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FADDX1_RVT S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FADDX1_RVT S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FADDX1_RVT S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), 
        .CO(\CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FADDX1_RVT S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), 
        .CO(\CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FADDX1_RVT S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), 
        .CO(\CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FADDX1_RVT S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), 
        .CO(\CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FADDX1_RVT S2_8_17 ( .A(\ab[8][17] ), .B(\CARRYB[7][17] ), .CI(\SUMB[7][18] ), .CO(\CARRYB[8][17] ), .S(\SUMB[8][17] ) );
  FADDX1_RVT S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), 
        .CO(\CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FADDX1_RVT S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), 
        .CO(\CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FADDX1_RVT S2_7_17 ( .A(\ab[7][17] ), .B(\CARRYB[6][17] ), .CI(\SUMB[6][18] ), .CO(\CARRYB[7][17] ), .S(\SUMB[7][17] ) );
  FADDX1_RVT S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), 
        .CO(\CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FADDX1_RVT S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), 
        .CO(\CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FADDX1_RVT S2_6_17 ( .A(\ab[6][17] ), .B(\CARRYB[5][17] ), .CI(\SUMB[5][18] ), .CO(\CARRYB[6][17] ), .S(\SUMB[6][17] ) );
  FADDX1_RVT S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), 
        .CO(\CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FADDX1_RVT S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), 
        .CO(\CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FADDX1_RVT S2_5_17 ( .A(\ab[5][17] ), .B(\CARRYB[4][17] ), .CI(\SUMB[4][18] ), .CO(\CARRYB[5][17] ), .S(\SUMB[5][17] ) );
  FADDX1_RVT S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), 
        .CO(\CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FADDX1_RVT S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), 
        .CO(\CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FADDX1_RVT S2_4_17 ( .A(\ab[4][17] ), .B(\CARRYB[3][17] ), .CI(\SUMB[3][18] ), .CO(\CARRYB[4][17] ), .S(\SUMB[4][17] ) );
  FADDX1_RVT S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), 
        .CO(\CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FADDX1_RVT S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), 
        .CO(\CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FADDX1_RVT S2_3_17 ( .A(\ab[3][17] ), .B(\CARRYB[2][17] ), .CI(\SUMB[2][18] ), .CO(\CARRYB[3][17] ), .S(\SUMB[3][17] ) );
  FADDX1_RVT S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), 
        .CO(\CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FADDX1_RVT S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), 
        .CO(\CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FADDX1_RVT S2_22_14 ( .A(\ab[22][14] ), .B(\CARRYB[21][14] ), .CI(
        \SUMB[21][15] ), .CO(\CARRYB[22][14] ), .S(\SUMB[22][14] ) );
  FADDX1_RVT S2_22_13 ( .A(\ab[22][13] ), .B(\CARRYB[21][13] ), .CI(
        \SUMB[21][14] ), .CO(\CARRYB[22][13] ), .S(\SUMB[22][13] ) );
  FADDX1_RVT S2_21_14 ( .A(\ab[21][14] ), .B(\CARRYB[20][14] ), .CI(
        \SUMB[20][15] ), .CO(\CARRYB[21][14] ), .S(\SUMB[21][14] ) );
  FADDX1_RVT S2_21_13 ( .A(\ab[21][13] ), .B(\CARRYB[20][13] ), .CI(
        \SUMB[20][14] ), .CO(\CARRYB[21][13] ), .S(\SUMB[21][13] ) );
  FADDX1_RVT S2_20_14 ( .A(\ab[20][14] ), .B(\CARRYB[19][14] ), .CI(
        \SUMB[19][15] ), .CO(\CARRYB[20][14] ), .S(\SUMB[20][14] ) );
  FADDX1_RVT S2_20_13 ( .A(\ab[20][13] ), .B(\CARRYB[19][13] ), .CI(
        \SUMB[19][14] ), .CO(\CARRYB[20][13] ), .S(\SUMB[20][13] ) );
  FADDX1_RVT S2_19_14 ( .A(\ab[19][14] ), .B(\CARRYB[18][14] ), .CI(
        \SUMB[18][15] ), .CO(\CARRYB[19][14] ), .S(\SUMB[19][14] ) );
  FADDX1_RVT S2_19_13 ( .A(\ab[19][13] ), .B(\CARRYB[18][13] ), .CI(
        \SUMB[18][14] ), .CO(\CARRYB[19][13] ), .S(\SUMB[19][13] ) );
  FADDX1_RVT S2_18_14 ( .A(\ab[18][14] ), .B(\CARRYB[17][14] ), .CI(
        \SUMB[17][15] ), .CO(\CARRYB[18][14] ), .S(\SUMB[18][14] ) );
  FADDX1_RVT S2_18_13 ( .A(\ab[18][13] ), .B(\CARRYB[17][13] ), .CI(
        \SUMB[17][14] ), .CO(\CARRYB[18][13] ), .S(\SUMB[18][13] ) );
  FADDX1_RVT S2_17_14 ( .A(\ab[17][14] ), .B(\CARRYB[16][14] ), .CI(
        \SUMB[16][15] ), .CO(\CARRYB[17][14] ), .S(\SUMB[17][14] ) );
  FADDX1_RVT S2_17_13 ( .A(\ab[17][13] ), .B(\CARRYB[16][13] ), .CI(
        \SUMB[16][14] ), .CO(\CARRYB[17][13] ), .S(\SUMB[17][13] ) );
  FADDX1_RVT S2_16_14 ( .A(\ab[16][14] ), .B(\CARRYB[15][14] ), .CI(
        \SUMB[15][15] ), .CO(\CARRYB[16][14] ), .S(\SUMB[16][14] ) );
  FADDX1_RVT S2_16_13 ( .A(\ab[16][13] ), .B(\CARRYB[15][13] ), .CI(
        \SUMB[15][14] ), .CO(\CARRYB[16][13] ), .S(\SUMB[16][13] ) );
  FADDX1_RVT S2_15_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(
        \SUMB[14][14] ), .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FADDX1_RVT S2_15_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(
        \SUMB[14][15] ), .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FADDX1_RVT S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(
        \SUMB[13][14] ), .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FADDX1_RVT S2_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(
        \SUMB[13][15] ), .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FADDX1_RVT S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(
        \SUMB[12][14] ), .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FADDX1_RVT S2_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(
        \SUMB[12][15] ), .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FADDX1_RVT S2_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(
        \SUMB[11][15] ), .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FADDX1_RVT S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(
        \SUMB[11][14] ), .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FADDX1_RVT S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(
        \SUMB[9][14] ), .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FADDX1_RVT S2_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(
        \SUMB[9][15] ), .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FADDX1_RVT S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FADDX1_RVT S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FADDX1_RVT S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FADDX1_RVT S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FADDX1_RVT S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FADDX1_RVT S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FADDX1_RVT S2_2_13 ( .A(\ab[2][13] ), .B(\CARRYB[1][13] ), .CI(\SUMB[1][14] ), .CO(\CARRYB[2][13] ), .S(\SUMB[2][13] ) );
  FADDX1_RVT S2_22_9 ( .A(\ab[22][9] ), .B(\CARRYB[21][9] ), .CI(
        \SUMB[21][10] ), .CO(\CARRYB[22][9] ), .S(\SUMB[22][9] ) );
  FADDX1_RVT S2_21_9 ( .A(\ab[21][9] ), .B(\CARRYB[20][9] ), .CI(
        \SUMB[20][10] ), .CO(\CARRYB[21][9] ), .S(\SUMB[21][9] ) );
  FADDX1_RVT S2_20_9 ( .A(\ab[20][9] ), .B(\CARRYB[19][9] ), .CI(
        \SUMB[19][10] ), .CO(\CARRYB[20][9] ), .S(\SUMB[20][9] ) );
  FADDX1_RVT S2_19_9 ( .A(\ab[19][9] ), .B(\CARRYB[18][9] ), .CI(
        \SUMB[18][10] ), .CO(\CARRYB[19][9] ), .S(\SUMB[19][9] ) );
  FADDX1_RVT S2_18_9 ( .A(\ab[18][9] ), .B(\CARRYB[17][9] ), .CI(
        \SUMB[17][10] ), .CO(\CARRYB[18][9] ), .S(\SUMB[18][9] ) );
  FADDX1_RVT S2_17_9 ( .A(\ab[17][9] ), .B(\CARRYB[16][9] ), .CI(
        \SUMB[16][10] ), .CO(\CARRYB[17][9] ), .S(\SUMB[17][9] ) );
  FADDX1_RVT S2_16_9 ( .A(\ab[16][9] ), .B(\CARRYB[15][9] ), .CI(
        \SUMB[15][10] ), .CO(\CARRYB[16][9] ), .S(\SUMB[16][9] ) );
  FADDX1_RVT S2_15_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(
        \SUMB[14][10] ), .CO(\CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FADDX1_RVT S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(
        \SUMB[13][10] ), .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FADDX1_RVT S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(
        \SUMB[12][10] ), .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FADDX1_RVT S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(
        \SUMB[11][10] ), .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FADDX1_RVT S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), 
        .CO(\CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FADDX1_RVT S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), 
        .CO(\CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FADDX1_RVT S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), 
        .CO(\CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FADDX1_RVT S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), 
        .CO(\CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FADDX1_RVT S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), 
        .CO(\CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FADDX1_RVT S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), 
        .CO(\CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FADDX1_RVT S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), 
        .CO(\CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FADDX1_RVT S2_2_9 ( .A(\ab[2][9] ), .B(\CARRYB[1][9] ), .CI(\SUMB[1][10] ), 
        .CO(\CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FADDX1_RVT S2_21_18 ( .A(\ab[21][18] ), .B(\CARRYB[20][18] ), .CI(
        \SUMB[20][19] ), .CO(\CARRYB[21][18] ), .S(\SUMB[21][18] ) );
  FADDX1_RVT S2_20_18 ( .A(\ab[20][18] ), .B(\CARRYB[19][18] ), .CI(
        \SUMB[19][19] ), .CO(\CARRYB[20][18] ), .S(\SUMB[20][18] ) );
  FADDX1_RVT S2_19_18 ( .A(\ab[19][18] ), .B(\CARRYB[18][18] ), .CI(
        \SUMB[18][19] ), .CO(\CARRYB[19][18] ), .S(\SUMB[19][18] ) );
  FADDX1_RVT S2_18_18 ( .A(\ab[18][18] ), .B(\CARRYB[17][18] ), .CI(
        \SUMB[17][19] ), .CO(\CARRYB[18][18] ), .S(\SUMB[18][18] ) );
  FADDX1_RVT S2_17_18 ( .A(\ab[17][18] ), .B(\CARRYB[16][18] ), .CI(
        \SUMB[16][19] ), .CO(\CARRYB[17][18] ), .S(\SUMB[17][18] ) );
  FADDX1_RVT S2_16_18 ( .A(\ab[16][18] ), .B(\CARRYB[15][18] ), .CI(
        \SUMB[15][19] ), .CO(\CARRYB[16][18] ), .S(\SUMB[16][18] ) );
  FADDX1_RVT S2_15_18 ( .A(\ab[15][18] ), .B(\CARRYB[14][18] ), .CI(
        \SUMB[14][19] ), .CO(\CARRYB[15][18] ), .S(\SUMB[15][18] ) );
  FADDX1_RVT S2_14_18 ( .A(\ab[14][18] ), .B(\CARRYB[13][18] ), .CI(
        \SUMB[13][19] ), .CO(\CARRYB[14][18] ), .S(\SUMB[14][18] ) );
  FADDX1_RVT S2_13_18 ( .A(\ab[13][18] ), .B(\CARRYB[12][18] ), .CI(
        \SUMB[12][19] ), .CO(\CARRYB[13][18] ), .S(\SUMB[13][18] ) );
  FADDX1_RVT S2_12_18 ( .A(\ab[12][18] ), .B(\CARRYB[11][18] ), .CI(
        \SUMB[11][19] ), .CO(\CARRYB[12][18] ), .S(\SUMB[12][18] ) );
  FADDX1_RVT S2_10_18 ( .A(\ab[10][18] ), .B(\CARRYB[9][18] ), .CI(
        \SUMB[9][19] ), .CO(\CARRYB[10][18] ), .S(\SUMB[10][18] ) );
  FADDX1_RVT S2_8_18 ( .A(\ab[8][18] ), .B(\CARRYB[7][18] ), .CI(\SUMB[7][19] ), .CO(\CARRYB[8][18] ), .S(\SUMB[8][18] ) );
  FADDX1_RVT S2_7_18 ( .A(\ab[7][18] ), .B(\CARRYB[6][18] ), .CI(\SUMB[6][19] ), .CO(\CARRYB[7][18] ), .S(\SUMB[7][18] ) );
  FADDX1_RVT S2_6_18 ( .A(\ab[6][18] ), .B(\CARRYB[5][18] ), .CI(\SUMB[5][19] ), .CO(\CARRYB[6][18] ), .S(\SUMB[6][18] ) );
  FADDX1_RVT S2_5_18 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .CI(\SUMB[4][19] ), .CO(\CARRYB[5][18] ), .S(\SUMB[5][18] ) );
  FADDX1_RVT S2_22_10 ( .A(\ab[22][10] ), .B(\CARRYB[21][10] ), .CI(
        \SUMB[21][11] ), .CO(\CARRYB[22][10] ), .S(\SUMB[22][10] ) );
  FADDX1_RVT S2_21_10 ( .A(\ab[21][10] ), .B(\CARRYB[20][10] ), .CI(
        \SUMB[20][11] ), .CO(\CARRYB[21][10] ), .S(\SUMB[21][10] ) );
  FADDX1_RVT S2_20_10 ( .A(\ab[20][10] ), .B(\CARRYB[19][10] ), .CI(
        \SUMB[19][11] ), .CO(\CARRYB[20][10] ), .S(\SUMB[20][10] ) );
  FADDX1_RVT S2_19_10 ( .A(\ab[19][10] ), .B(\CARRYB[18][10] ), .CI(
        \SUMB[18][11] ), .CO(\CARRYB[19][10] ), .S(\SUMB[19][10] ) );
  FADDX1_RVT S2_18_10 ( .A(\ab[18][10] ), .B(\CARRYB[17][10] ), .CI(
        \SUMB[17][11] ), .CO(\CARRYB[18][10] ), .S(\SUMB[18][10] ) );
  FADDX1_RVT S2_17_10 ( .A(\ab[17][10] ), .B(\CARRYB[16][10] ), .CI(
        \SUMB[16][11] ), .CO(\CARRYB[17][10] ), .S(\SUMB[17][10] ) );
  FADDX1_RVT S2_16_10 ( .A(\ab[16][10] ), .B(\CARRYB[15][10] ), .CI(
        \SUMB[15][11] ), .CO(\CARRYB[16][10] ), .S(\SUMB[16][10] ) );
  FADDX1_RVT S2_15_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(
        \SUMB[14][11] ), .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FADDX1_RVT S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(
        \SUMB[13][11] ), .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FADDX1_RVT S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(
        \SUMB[12][11] ), .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FADDX1_RVT S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(
        \SUMB[9][11] ), .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FADDX1_RVT S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FADDX1_RVT S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FADDX1_RVT S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FADDX1_RVT S2_22_5 ( .A(\ab[22][5] ), .B(\CARRYB[21][5] ), .CI(\SUMB[21][6] ), .CO(\CARRYB[22][5] ), .S(\SUMB[22][5] ) );
  FADDX1_RVT S2_21_5 ( .A(\ab[21][5] ), .B(\CARRYB[20][5] ), .CI(\SUMB[20][6] ), .CO(\CARRYB[21][5] ), .S(\SUMB[21][5] ) );
  FADDX1_RVT S2_20_5 ( .A(\ab[20][5] ), .B(\CARRYB[19][5] ), .CI(\SUMB[19][6] ), .CO(\CARRYB[20][5] ), .S(\SUMB[20][5] ) );
  FADDX1_RVT S2_19_5 ( .A(\ab[19][5] ), .B(\CARRYB[18][5] ), .CI(\SUMB[18][6] ), .CO(\CARRYB[19][5] ), .S(\SUMB[19][5] ) );
  FADDX1_RVT S2_18_5 ( .A(\ab[18][5] ), .B(\CARRYB[17][5] ), .CI(\SUMB[17][6] ), .CO(\CARRYB[18][5] ), .S(\SUMB[18][5] ) );
  FADDX1_RVT S2_17_5 ( .A(\ab[17][5] ), .B(\CARRYB[16][5] ), .CI(\SUMB[16][6] ), .CO(\CARRYB[17][5] ), .S(\SUMB[17][5] ) );
  FADDX1_RVT S2_16_5 ( .A(\ab[16][5] ), .B(\CARRYB[15][5] ), .CI(\SUMB[15][6] ), .CO(\CARRYB[16][5] ), .S(\SUMB[16][5] ) );
  FADDX1_RVT S2_15_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), .CO(\CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FADDX1_RVT S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FADDX1_RVT S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FADDX1_RVT S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FADDX1_RVT S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), 
        .CO(\CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FADDX1_RVT S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), 
        .CO(\CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FADDX1_RVT S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), 
        .CO(\CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FADDX1_RVT S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), 
        .CO(\CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FADDX1_RVT S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), 
        .CO(\CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FADDX1_RVT S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), 
        .CO(\CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FADDX1_RVT S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), 
        .CO(\CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FADDX1_RVT S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), 
        .CO(\CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FADDX1_RVT S2_3_21 ( .A(\ab[3][21] ), .B(\CARRYB[2][21] ), .CI(\SUMB[2][22] ), .CO(\CARRYB[3][21] ), .S(\SUMB[3][21] ) );
  FADDX1_RVT S2_22_15 ( .A(\ab[22][15] ), .B(\CARRYB[21][15] ), .CI(
        \SUMB[21][16] ), .CO(\CARRYB[22][15] ), .S(\SUMB[22][15] ) );
  FADDX1_RVT S2_21_15 ( .A(\ab[21][15] ), .B(\CARRYB[20][15] ), .CI(
        \SUMB[20][16] ), .CO(\CARRYB[21][15] ), .S(\SUMB[21][15] ) );
  FADDX1_RVT S2_20_15 ( .A(\ab[20][15] ), .B(\CARRYB[19][15] ), .CI(
        \SUMB[19][16] ), .CO(\CARRYB[20][15] ), .S(\SUMB[20][15] ) );
  FADDX1_RVT S2_22_11 ( .A(\ab[22][11] ), .B(\CARRYB[21][11] ), .CI(
        \SUMB[21][12] ), .CO(\CARRYB[22][11] ), .S(\SUMB[22][11] ) );
  FADDX1_RVT S2_19_15 ( .A(\ab[19][15] ), .B(\CARRYB[18][15] ), .CI(
        \SUMB[18][16] ), .CO(\CARRYB[19][15] ), .S(\SUMB[19][15] ) );
  FADDX1_RVT S2_21_11 ( .A(\ab[21][11] ), .B(\CARRYB[20][11] ), .CI(
        \SUMB[20][12] ), .CO(\CARRYB[21][11] ), .S(\SUMB[21][11] ) );
  FADDX1_RVT S2_18_15 ( .A(\ab[18][15] ), .B(\CARRYB[17][15] ), .CI(
        \SUMB[17][16] ), .CO(\CARRYB[18][15] ), .S(\SUMB[18][15] ) );
  FADDX1_RVT S2_20_11 ( .A(\ab[20][11] ), .B(\CARRYB[19][11] ), .CI(
        \SUMB[19][12] ), .CO(\CARRYB[20][11] ), .S(\SUMB[20][11] ) );
  FADDX1_RVT S2_17_15 ( .A(\ab[17][15] ), .B(\CARRYB[16][15] ), .CI(
        \SUMB[16][16] ), .CO(\CARRYB[17][15] ), .S(\SUMB[17][15] ) );
  FADDX1_RVT S2_19_11 ( .A(\ab[19][11] ), .B(\CARRYB[18][11] ), .CI(
        \SUMB[18][12] ), .CO(\CARRYB[19][11] ), .S(\SUMB[19][11] ) );
  FADDX1_RVT S2_16_15 ( .A(\ab[16][15] ), .B(\CARRYB[15][15] ), .CI(
        \SUMB[15][16] ), .CO(\CARRYB[16][15] ), .S(\SUMB[16][15] ) );
  FADDX1_RVT S2_18_11 ( .A(\ab[18][11] ), .B(\CARRYB[17][11] ), .CI(
        \SUMB[17][12] ), .CO(\CARRYB[18][11] ), .S(\SUMB[18][11] ) );
  FADDX1_RVT S2_17_11 ( .A(\ab[17][11] ), .B(\CARRYB[16][11] ), .CI(
        \SUMB[16][12] ), .CO(\CARRYB[17][11] ), .S(\SUMB[17][11] ) );
  FADDX1_RVT S2_15_15 ( .A(\ab[15][15] ), .B(\CARRYB[14][15] ), .CI(
        \SUMB[14][16] ), .CO(\CARRYB[15][15] ), .S(\SUMB[15][15] ) );
  FADDX1_RVT S2_16_11 ( .A(\ab[16][11] ), .B(\CARRYB[15][11] ), .CI(
        \SUMB[15][12] ), .CO(\CARRYB[16][11] ), .S(\SUMB[16][11] ) );
  FADDX1_RVT S2_15_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(
        \SUMB[14][12] ), .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FADDX1_RVT S2_14_15 ( .A(\ab[14][15] ), .B(\CARRYB[13][15] ), .CI(
        \SUMB[13][16] ), .CO(\CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FADDX1_RVT S2_13_15 ( .A(\ab[13][15] ), .B(\CARRYB[12][15] ), .CI(
        \SUMB[12][16] ), .CO(\CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FADDX1_RVT S2_12_15 ( .A(\ab[12][15] ), .B(\CARRYB[11][15] ), .CI(
        \SUMB[11][16] ), .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FADDX1_RVT S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(
        \SUMB[13][12] ), .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FADDX1_RVT S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(
        \SUMB[12][12] ), .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FADDX1_RVT S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(
        \SUMB[11][12] ), .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FADDX1_RVT S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(
        \SUMB[9][12] ), .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FADDX1_RVT S2_10_15 ( .A(\ab[10][15] ), .B(\CARRYB[9][15] ), .CI(
        \SUMB[9][16] ), .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FADDX1_RVT S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FADDX1_RVT S2_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\SUMB[7][16] ), .CO(\CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FADDX1_RVT S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FADDX1_RVT S2_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\SUMB[6][16] ), .CO(\CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FADDX1_RVT S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FADDX1_RVT S2_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .CI(\SUMB[5][16] ), .CO(\CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FADDX1_RVT S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FADDX1_RVT S2_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .CI(\SUMB[4][16] ), .CO(\CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FADDX1_RVT S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FADDX1_RVT S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\SUMB[3][16] ), .CO(\CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FADDX1_RVT S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FADDX1_RVT S2_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .CI(\SUMB[2][16] ), .CO(\CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FADDX1_RVT S2_2_11 ( .A(\ab[2][11] ), .B(\CARRYB[1][11] ), .CI(\SUMB[1][12] ), .CO(\CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FADDX1_RVT S2_2_15 ( .A(\ab[2][15] ), .B(\CARRYB[1][15] ), .CI(\SUMB[1][16] ), .CO(\CARRYB[2][15] ), .S(\SUMB[2][15] ) );
  FADDX1_RVT S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), 
        .CO(\CARRYB[9][0] ), .S(\A1[7] ) );
  FADDX1_RVT S2_20_19 ( .A(\ab[20][19] ), .B(\CARRYB[19][19] ), .CI(
        \SUMB[19][20] ), .CO(\CARRYB[20][19] ), .S(\SUMB[20][19] ) );
  FADDX1_RVT S2_19_19 ( .A(\ab[19][19] ), .B(\CARRYB[18][19] ), .CI(
        \SUMB[18][20] ), .CO(\CARRYB[19][19] ), .S(\SUMB[19][19] ) );
  FADDX1_RVT S2_18_19 ( .A(\ab[18][19] ), .B(\CARRYB[17][19] ), .CI(
        \SUMB[17][20] ), .CO(\CARRYB[18][19] ), .S(\SUMB[18][19] ) );
  FADDX1_RVT S2_17_19 ( .A(\ab[17][19] ), .B(\CARRYB[16][19] ), .CI(
        \SUMB[16][20] ), .CO(\CARRYB[17][19] ), .S(\SUMB[17][19] ) );
  FADDX1_RVT S2_16_19 ( .A(\ab[16][19] ), .B(\CARRYB[15][19] ), .CI(
        \SUMB[15][20] ), .CO(\CARRYB[16][19] ), .S(\SUMB[16][19] ) );
  FADDX1_RVT S2_15_19 ( .A(\ab[15][19] ), .B(\CARRYB[14][19] ), .CI(
        \SUMB[14][20] ), .CO(\CARRYB[15][19] ), .S(\SUMB[15][19] ) );
  FADDX1_RVT S2_14_19 ( .A(\ab[14][19] ), .B(\CARRYB[13][19] ), .CI(
        \SUMB[13][20] ), .CO(\CARRYB[14][19] ), .S(\SUMB[14][19] ) );
  FADDX1_RVT S2_13_19 ( .A(\ab[13][19] ), .B(\CARRYB[12][19] ), .CI(
        \SUMB[12][20] ), .CO(\CARRYB[13][19] ), .S(\SUMB[13][19] ) );
  FADDX1_RVT S2_12_19 ( .A(\ab[12][19] ), .B(\CARRYB[11][19] ), .CI(
        \SUMB[11][20] ), .CO(\CARRYB[12][19] ), .S(\SUMB[12][19] ) );
  FADDX1_RVT S2_10_19 ( .A(\ab[10][19] ), .B(\CARRYB[9][19] ), .CI(
        \SUMB[9][20] ), .CO(\CARRYB[10][19] ), .S(\SUMB[10][19] ) );
  FADDX1_RVT S2_8_19 ( .A(\ab[8][19] ), .B(\CARRYB[7][19] ), .CI(\SUMB[7][20] ), .CO(\CARRYB[8][19] ), .S(\SUMB[8][19] ) );
  FADDX1_RVT S2_7_19 ( .A(\ab[7][19] ), .B(\CARRYB[6][19] ), .CI(\SUMB[6][20] ), .CO(\CARRYB[7][19] ), .S(\SUMB[7][19] ) );
  FADDX1_RVT S2_6_19 ( .A(\ab[6][19] ), .B(\CARRYB[5][19] ), .CI(\SUMB[5][20] ), .CO(\CARRYB[6][19] ), .S(\SUMB[6][19] ) );
  FADDX1_RVT S2_5_19 ( .A(\ab[5][19] ), .B(\CARRYB[4][19] ), .CI(\SUMB[4][20] ), .CO(\CARRYB[5][19] ), .S(\SUMB[5][19] ) );
  FADDX1_RVT S2_4_19 ( .A(\ab[4][19] ), .B(\CARRYB[3][19] ), .CI(\SUMB[3][20] ), .CO(\CARRYB[4][19] ), .S(\SUMB[4][19] ) );
  FADDX1_RVT S2_3_19 ( .A(\ab[3][19] ), .B(\CARRYB[2][19] ), .CI(\SUMB[2][20] ), .CO(\CARRYB[3][19] ), .S(\SUMB[3][19] ) );
  FADDX1_RVT S2_2_19 ( .A(\ab[2][19] ), .B(\CARRYB[1][19] ), .CI(\SUMB[1][20] ), .CO(\CARRYB[2][19] ), .S(\SUMB[2][19] ) );
  FADDX1_RVT S2_12_21 ( .A(\ab[12][21] ), .B(\CARRYB[11][21] ), .CI(
        \SUMB[11][22] ), .CO(\CARRYB[12][21] ), .S(\SUMB[12][21] ) );
  FADDX1_RVT S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), 
        .CO(\CARRYB[6][0] ), .S(\A1[4] ) );
  FADDX1_RVT S1_16_0 ( .A(\ab[16][0] ), .B(\CARRYB[15][0] ), .CI(\SUMB[15][1] ), .CO(\CARRYB[16][0] ), .S(\A1[14] ) );
  FADDX1_RVT S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FADDX1_RVT S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), 
        .CO(\CARRYB[4][0] ), .S(\A1[2] ) );
  FADDX1_RVT S1_17_0 ( .A(\ab[17][0] ), .B(\CARRYB[16][0] ), .CI(\SUMB[16][1] ), .CO(\CARRYB[17][0] ), .S(\A1[15] ) );
  FADDX1_RVT S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), 
        .CO(\CARRYB[7][0] ), .S(\A1[5] ) );
  FADDX1_RVT S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FADDX1_RVT S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), .CO(\CARRYB[14][0] ), .S(\A1[12] ) );
  FADDX1_RVT S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), 
        .CO(\CARRYB[3][0] ), .S(\A1[1] ) );
  FADDX1_RVT S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), 
        .CO(\CARRYB[8][0] ), .S(\A1[6] ) );
  FADDX1_RVT S1_20_0 ( .A(\ab[20][0] ), .B(\CARRYB[19][0] ), .CI(\SUMB[19][1] ), .CO(\CARRYB[20][0] ), .S(\A1[18] ) );
  FADDX1_RVT S1_18_0 ( .A(\ab[18][0] ), .B(\CARRYB[17][0] ), .CI(\SUMB[17][1] ), .CO(\CARRYB[18][0] ), .S(\A1[16] ) );
  FADDX1_RVT S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), 
        .CO(\CARRYB[5][0] ), .S(\A1[3] ) );
  FADDX1_RVT S1_15_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), .CO(\CARRYB[15][0] ), .S(\A1[13] ) );
  FADDX1_RVT S2_20_2 ( .A(\ab[20][2] ), .B(\CARRYB[19][2] ), .CI(\SUMB[19][3] ), .CO(\CARRYB[20][2] ), .S(\SUMB[20][2] ) );
  FADDX1_RVT S2_18_2 ( .A(\ab[18][2] ), .B(\CARRYB[17][2] ), .CI(\SUMB[17][3] ), .CO(\CARRYB[18][2] ), .S(\SUMB[18][2] ) );
  FADDX1_RVT S2_17_2 ( .A(\ab[17][2] ), .B(\CARRYB[16][2] ), .CI(\SUMB[16][3] ), .CO(\CARRYB[17][2] ), .S(\SUMB[17][2] ) );
  FADDX1_RVT S2_16_2 ( .A(\ab[16][2] ), .B(\CARRYB[15][2] ), .CI(\SUMB[15][3] ), .CO(\CARRYB[16][2] ), .S(\SUMB[16][2] ) );
  FADDX1_RVT S2_15_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), .CO(\CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FADDX1_RVT S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FADDX1_RVT S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FADDX1_RVT S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FADDX1_RVT S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), 
        .CO(\CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FADDX1_RVT S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), 
        .CO(\CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FADDX1_RVT S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), 
        .CO(\CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FADDX1_RVT S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), 
        .CO(\CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FADDX1_RVT S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), 
        .CO(\CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FADDX1_RVT S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), 
        .CO(\CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FADDX1_RVT S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), 
        .CO(\CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FADDX1_RVT S1_19_0 ( .A(\ab[19][0] ), .B(\CARRYB[18][0] ), .CI(\SUMB[18][1] ), .CO(\CARRYB[19][0] ), .S(\A1[17] ) );
  FADDX1_RVT S2_19_2 ( .A(\ab[19][2] ), .B(\CARRYB[18][2] ), .CI(\SUMB[18][3] ), .CO(\CARRYB[19][2] ), .S(\SUMB[19][2] ) );
  FADDX1_RVT S2_4_21 ( .A(\ab[4][21] ), .B(\CARRYB[3][21] ), .CI(\SUMB[3][22] ), .CO(\CARRYB[4][21] ), .S(\SUMB[4][21] ) );
  FADDX1_RVT S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FADDX1_RVT S2_11_20 ( .A(\ab[11][20] ), .B(\CARRYB[10][20] ), .CI(
        \SUMB[10][21] ), .CO(\CARRYB[11][20] ), .S(\SUMB[11][20] ) );
  FADDX1_RVT S2_11_19 ( .A(\ab[11][19] ), .B(\CARRYB[10][19] ), .CI(
        \SUMB[10][20] ), .CO(\CARRYB[11][19] ), .S(\SUMB[11][19] ) );
  FADDX1_RVT S2_11_15 ( .A(\ab[11][15] ), .B(\CARRYB[10][15] ), .CI(
        \SUMB[10][16] ), .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FADDX1_RVT S2_11_16 ( .A(\ab[11][16] ), .B(\CARRYB[10][16] ), .CI(
        \SUMB[10][17] ), .CO(\CARRYB[11][16] ), .S(\SUMB[11][16] ) );
  FADDX1_RVT S2_11_17 ( .A(\ab[11][17] ), .B(\CARRYB[10][17] ), .CI(
        \SUMB[10][18] ), .CO(\CARRYB[11][17] ), .S(\SUMB[11][17] ) );
  FADDX1_RVT S2_11_18 ( .A(\ab[11][18] ), .B(\CARRYB[10][18] ), .CI(
        \SUMB[10][19] ), .CO(\CARRYB[11][18] ), .S(\SUMB[11][18] ) );
  FADDX1_RVT S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FADDX1_RVT S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FADDX1_RVT S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FADDX1_RVT S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FADDX1_RVT S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FADDX1_RVT S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FADDX1_RVT S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(
        \SUMB[10][10] ), .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FADDX1_RVT S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(
        \SUMB[10][11] ), .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FADDX1_RVT S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(
        \SUMB[10][12] ), .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FADDX1_RVT S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(
        \SUMB[10][13] ), .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FADDX1_RVT S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(
        \SUMB[10][14] ), .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FADDX1_RVT S2_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(
        \SUMB[10][15] ), .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FADDX1_RVT S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), 
        .CO(\CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FADDX1_RVT S2_9_16 ( .A(\ab[9][16] ), .B(\CARRYB[8][16] ), .CI(\SUMB[8][17] ), .CO(\CARRYB[9][16] ), .S(\SUMB[9][16] ) );
  FADDX1_RVT S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FADDX1_RVT S2_9_20 ( .A(\ab[9][20] ), .B(\CARRYB[8][20] ), .CI(\SUMB[8][21] ), .CO(\CARRYB[9][20] ), .S(\SUMB[9][20] ) );
  FADDX1_RVT S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), 
        .CO(\CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FADDX1_RVT S2_9_17 ( .A(\ab[9][17] ), .B(\CARRYB[8][17] ), .CI(\SUMB[8][18] ), .CO(\CARRYB[9][17] ), .S(\SUMB[9][17] ) );
  FADDX1_RVT S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), 
        .CO(\CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FADDX1_RVT S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), 
        .CO(\CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FADDX1_RVT S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FADDX1_RVT S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FADDX1_RVT S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), 
        .CO(\CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FADDX1_RVT S2_9_18 ( .A(\ab[9][18] ), .B(\CARRYB[8][18] ), .CI(\SUMB[8][19] ), .CO(\CARRYB[9][18] ), .S(\SUMB[9][18] ) );
  FADDX1_RVT S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FADDX1_RVT S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), 
        .CO(\CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FADDX1_RVT S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(
        \SUMB[9][13] ), .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FADDX1_RVT S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FADDX1_RVT S2_9_15 ( .A(\ab[9][15] ), .B(\CARRYB[8][15] ), .CI(\SUMB[8][16] ), .CO(\CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FADDX1_RVT S2_18_4 ( .A(\ab[18][4] ), .B(\CARRYB[17][4] ), .CI(\SUMB[17][5] ), .CO(\CARRYB[18][4] ), .S(\SUMB[18][4] ) );
  FADDX1_RVT S2_17_4 ( .A(\ab[17][4] ), .B(\CARRYB[16][4] ), .CI(\SUMB[16][5] ), .CO(\CARRYB[17][4] ), .S(\SUMB[17][4] ) );
  FADDX1_RVT S2_16_4 ( .A(\ab[16][4] ), .B(\CARRYB[15][4] ), .CI(\SUMB[15][5] ), .CO(\CARRYB[16][4] ), .S(\SUMB[16][4] ) );
  FADDX1_RVT S2_15_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), .CO(\CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FADDX1_RVT S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FADDX1_RVT S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FADDX1_RVT S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FADDX1_RVT S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FADDX1_RVT S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), 
        .CO(\CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FADDX1_RVT S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), 
        .CO(\CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FADDX1_RVT S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), 
        .CO(\CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FADDX1_RVT S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), 
        .CO(\CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FADDX1_RVT S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), 
        .CO(\CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FADDX1_RVT S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), 
        .CO(\CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FADDX1_RVT S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), 
        .CO(\CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FADDX1_RVT S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), 
        .CO(\CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FADDX1_RVT S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), 
        .CO(\CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FADDX1_RVT S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), 
        .CO(\CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FADDX1_RVT S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), 
        .CO(\CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FADDX1_RVT S2_2_8 ( .A(\ab[2][8] ), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), 
        .CO(\CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FADDX1_RVT S2_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FADDX1_RVT S2_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FADDX1_RVT S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\SUMB[5][15] ), .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FADDX1_RVT S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FADDX1_RVT S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FADDX1_RVT S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FADDX1_RVT S2_2_14 ( .A(\ab[2][14] ), .B(\CARRYB[1][14] ), .CI(\SUMB[1][15] ), .CO(\CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  FADDX1_RVT S2_9_19 ( .A(\ab[9][19] ), .B(\CARRYB[8][19] ), .CI(\SUMB[8][20] ), .CO(\CARRYB[9][19] ), .S(\SUMB[9][19] ) );
  FADDX1_RVT S2_4_18 ( .A(\ab[4][18] ), .B(\CARRYB[3][18] ), .CI(\SUMB[3][19] ), .CO(\CARRYB[4][18] ), .S(\SUMB[4][18] ) );
  FADDX1_RVT S2_3_18 ( .A(\ab[3][18] ), .B(\CARRYB[2][18] ), .CI(\SUMB[2][19] ), .CO(\CARRYB[3][18] ), .S(\SUMB[3][18] ) );
  FADDX1_RVT S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(
        \SUMB[11][11] ), .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FADDX1_RVT S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FADDX1_RVT S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FADDX1_RVT S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FADDX1_RVT S2_2_10 ( .A(\ab[2][10] ), .B(\CARRYB[1][10] ), .CI(\SUMB[1][11] ), .CO(\CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FADDX1_RVT S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), 
        .CO(\CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FADDX1_RVT S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FADDX1_RVT S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FADDX1_RVT S2_8_21 ( .A(\ab[8][21] ), .B(\CARRYB[7][21] ), .CI(\SUMB[7][22] ), .CO(\CARRYB[8][21] ), .S(\SUMB[8][21] ) );
  FADDX1_RVT S2_18_21 ( .A(\ab[18][21] ), .B(\CARRYB[17][21] ), .CI(
        \SUMB[17][22] ), .CO(\CARRYB[18][21] ), .S(\SUMB[18][21] ) );
  FADDX1_RVT S2_14_21 ( .A(\ab[14][21] ), .B(\CARRYB[13][21] ), .CI(
        \SUMB[13][22] ), .CO(\CARRYB[14][21] ), .S(\SUMB[14][21] ) );
  FADDX1_RVT S2_6_21 ( .A(\ab[6][21] ), .B(\CARRYB[5][21] ), .CI(\SUMB[5][22] ), .CO(\CARRYB[6][21] ), .S(\SUMB[6][21] ) );
  FADDX1_RVT S2_9_21 ( .A(\ab[9][21] ), .B(\CARRYB[8][21] ), .CI(\SUMB[8][22] ), .CO(\CARRYB[9][21] ), .S(\SUMB[9][21] ) );
  FADDX1_RVT S2_15_21 ( .A(\ab[15][21] ), .B(\CARRYB[14][21] ), .CI(
        \SUMB[14][22] ), .CO(\CARRYB[15][21] ), .S(\SUMB[15][21] ) );
  FADDX1_RVT S2_5_21 ( .A(\ab[5][21] ), .B(\CARRYB[4][21] ), .CI(\SUMB[4][22] ), .CO(\CARRYB[5][21] ), .S(\SUMB[5][21] ) );
  FADDX1_RVT S2_16_21 ( .A(\ab[16][21] ), .B(\CARRYB[15][21] ), .CI(
        \SUMB[15][22] ), .CO(\CARRYB[16][21] ), .S(\SUMB[16][21] ) );
  FADDX1_RVT S2_11_21 ( .A(\ab[11][21] ), .B(\CARRYB[10][21] ), .CI(
        \SUMB[10][22] ), .CO(\CARRYB[11][21] ), .S(\SUMB[11][21] ) );
  FADDX1_RVT S2_10_21 ( .A(\ab[10][21] ), .B(\CARRYB[9][21] ), .CI(
        \SUMB[9][22] ), .CO(\CARRYB[10][21] ), .S(\SUMB[10][21] ) );
  FADDX1_RVT S2_7_21 ( .A(\ab[7][21] ), .B(\CARRYB[6][21] ), .CI(\SUMB[6][22] ), .CO(\CARRYB[7][21] ), .S(\SUMB[7][21] ) );
  FADDX1_RVT S2_17_21 ( .A(\ab[17][21] ), .B(\CARRYB[16][21] ), .CI(
        \SUMB[16][22] ), .CO(\CARRYB[17][21] ), .S(\SUMB[17][21] ) );
  FADDX1_RVT S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), 
        .CO(\CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FADDX1_RVT S2_13_21 ( .A(\ab[13][21] ), .B(\CARRYB[12][21] ), .CI(
        \SUMB[12][22] ), .CO(\CARRYB[13][21] ), .S(\SUMB[13][21] ) );
  FADDX1_RVT S2_2_21 ( .A(\ab[2][21] ), .B(\CARRYB[1][21] ), .CI(\SUMB[1][22] ), .CO(\CARRYB[2][21] ), .S(\SUMB[2][21] ) );
  FADDX1_RVT S3_2_22 ( .A(\ab[2][22] ), .B(\CARRYB[1][22] ), .CI(n51), .CO(
        \CARRYB[2][22] ), .S(\SUMB[2][22] ) );
  FADDX1_RVT S4_1 ( .A(n5), .B(\CARRYB[22][1] ), .CI(\SUMB[22][2] ), .CO(
        \CARRYB[23][1] ), .S(\SUMB[23][1] ) );
  FADDX1_RVT S4_0 ( .A(n3), .B(\CARRYB[22][0] ), .CI(\SUMB[22][1] ), .CO(
        \CARRYB[23][0] ), .S(\SUMB[23][0] ) );
  FADDX1_RVT S3_11_22 ( .A(\ab[11][22] ), .B(\CARRYB[10][22] ), .CI(n69), .CO(
        \CARRYB[11][22] ), .S(\SUMB[11][22] ) );
  FADDX1_RVT S3_3_22 ( .A(\ab[3][22] ), .B(\CARRYB[2][22] ), .CI(n53), .CO(
        \CARRYB[3][22] ), .S(\SUMB[3][22] ) );
  FADDX1_RVT S4_2 ( .A(n7), .B(\CARRYB[22][2] ), .CI(\SUMB[22][3] ), .CO(
        \CARRYB[23][2] ), .S(\SUMB[23][2] ) );
  FADDX1_RVT S4_16 ( .A(n35), .B(\CARRYB[22][16] ), .CI(\SUMB[22][17] ), .CO(
        \CARRYB[23][16] ), .S(\SUMB[23][16] ) );
  FADDX1_RVT S4_6 ( .A(n15), .B(\CARRYB[22][6] ), .CI(\SUMB[22][7] ), .CO(
        \CARRYB[23][6] ), .S(\SUMB[23][6] ) );
  FADDX1_RVT S4_12 ( .A(n27), .B(\CARRYB[22][12] ), .CI(\SUMB[22][13] ), .CO(
        \CARRYB[23][12] ), .S(\SUMB[23][12] ) );
  FADDX1_RVT S4_4 ( .A(n11), .B(\CARRYB[22][4] ), .CI(\SUMB[22][5] ), .CO(
        \CARRYB[23][4] ), .S(\SUMB[23][4] ) );
  FADDX1_RVT S4_8 ( .A(n19), .B(\CARRYB[22][8] ), .CI(\SUMB[22][9] ), .CO(
        \CARRYB[23][8] ), .S(\SUMB[23][8] ) );
  FADDX1_RVT S4_3 ( .A(n9), .B(\CARRYB[22][3] ), .CI(\SUMB[22][4] ), .CO(
        \CARRYB[23][3] ), .S(\SUMB[23][3] ) );
  FADDX1_RVT S4_7 ( .A(n17), .B(\CARRYB[22][7] ), .CI(\SUMB[22][8] ), .CO(
        \CARRYB[23][7] ), .S(\SUMB[23][7] ) );
  FADDX1_RVT S4_14 ( .A(n31), .B(\CARRYB[22][14] ), .CI(\SUMB[22][15] ), .CO(
        \CARRYB[23][14] ), .S(\SUMB[23][14] ) );
  FADDX1_RVT S4_13 ( .A(n29), .B(\CARRYB[22][13] ), .CI(\SUMB[22][14] ), .CO(
        \CARRYB[23][13] ), .S(\SUMB[23][13] ) );
  FADDX1_RVT S4_9 ( .A(n21), .B(\CARRYB[22][9] ), .CI(\SUMB[22][10] ), .CO(
        \CARRYB[23][9] ), .S(\SUMB[23][9] ) );
  FADDX1_RVT S4_10 ( .A(n23), .B(\CARRYB[22][10] ), .CI(\SUMB[22][11] ), .CO(
        \CARRYB[23][10] ), .S(\SUMB[23][10] ) );
  FADDX1_RVT S4_5 ( .A(n13), .B(\CARRYB[22][5] ), .CI(\SUMB[22][6] ), .CO(
        \CARRYB[23][5] ), .S(\SUMB[23][5] ) );
  FADDX1_RVT S4_15 ( .A(n33), .B(\CARRYB[22][15] ), .CI(\SUMB[22][16] ), .CO(
        \CARRYB[23][15] ), .S(\SUMB[23][15] ) );
  FADDX1_RVT S4_11 ( .A(n25), .B(\CARRYB[22][11] ), .CI(\SUMB[22][12] ), .CO(
        \CARRYB[23][11] ), .S(\SUMB[23][11] ) );
  FADDX1_RVT S3_7_22 ( .A(\ab[7][22] ), .B(\CARRYB[6][22] ), .CI(n61), .CO(
        \CARRYB[7][22] ), .S(\SUMB[7][22] ) );
  FADDX1_RVT S3_17_22 ( .A(\ab[17][22] ), .B(\CARRYB[16][22] ), .CI(n81), .CO(
        \CARRYB[17][22] ), .S(\SUMB[17][22] ) );
  FADDX1_RVT S3_13_22 ( .A(\ab[13][22] ), .B(\CARRYB[12][22] ), .CI(n73), .CO(
        \CARRYB[13][22] ), .S(\SUMB[13][22] ) );
  FADDX1_RVT S3_5_22 ( .A(\ab[5][22] ), .B(\CARRYB[4][22] ), .CI(n57), .CO(
        \CARRYB[5][22] ), .S(\SUMB[5][22] ) );
  FADDX1_RVT S3_8_22 ( .A(\ab[8][22] ), .B(\CARRYB[7][22] ), .CI(n63), .CO(
        \CARRYB[8][22] ), .S(\SUMB[8][22] ) );
  FADDX1_RVT S3_14_22 ( .A(\ab[14][22] ), .B(\CARRYB[13][22] ), .CI(n75), .CO(
        \CARRYB[14][22] ), .S(\SUMB[14][22] ) );
  FADDX1_RVT S3_4_22 ( .A(\ab[4][22] ), .B(\CARRYB[3][22] ), .CI(n55), .CO(
        \CARRYB[4][22] ), .S(\SUMB[4][22] ) );
  FADDX1_RVT S3_15_22 ( .A(\ab[15][22] ), .B(\CARRYB[14][22] ), .CI(n77), .CO(
        \CARRYB[15][22] ), .S(\SUMB[15][22] ) );
  FADDX1_RVT S3_10_22 ( .A(\ab[10][22] ), .B(\CARRYB[9][22] ), .CI(n67), .CO(
        \CARRYB[10][22] ), .S(\SUMB[10][22] ) );
  FADDX1_RVT S3_9_22 ( .A(\ab[9][22] ), .B(\CARRYB[8][22] ), .CI(n65), .CO(
        \CARRYB[9][22] ), .S(\SUMB[9][22] ) );
  FADDX1_RVT S3_6_22 ( .A(\ab[6][22] ), .B(\CARRYB[5][22] ), .CI(n59), .CO(
        \CARRYB[6][22] ), .S(\SUMB[6][22] ) );
  FADDX1_RVT S3_16_22 ( .A(\ab[16][22] ), .B(\CARRYB[15][22] ), .CI(n79), .CO(
        \CARRYB[16][22] ), .S(\SUMB[16][22] ) );
  FADDX1_RVT S3_12_22 ( .A(\ab[12][22] ), .B(\CARRYB[11][22] ), .CI(n71), .CO(
        \CARRYB[12][22] ), .S(\SUMB[12][22] ) );
  INVX0_RVT U2 ( .A(\ab[5][23] ), .Y(n60) );
  INVX0_RVT U3 ( .A(\ab[4][23] ), .Y(n58) );
  INVX0_RVT U4 ( .A(\ab[20][23] ), .Y(n90) );
  INVX0_RVT U5 ( .A(\ab[16][23] ), .Y(n82) );
  INVX0_RVT U6 ( .A(\ab[13][23] ), .Y(n76) );
  INVX0_RVT U7 ( .A(\ab[18][23] ), .Y(n86) );
  INVX0_RVT U8 ( .A(\ab[15][23] ), .Y(n80) );
  INVX0_RVT U9 ( .A(\ab[12][23] ), .Y(n74) );
  INVX0_RVT U10 ( .A(\ab[17][23] ), .Y(n84) );
  INVX0_RVT U11 ( .A(\ab[11][23] ), .Y(n72) );
  INVX1_RVT U12 ( .A(n58), .Y(n57) );
  INVX1_RVT U13 ( .A(n74), .Y(n73) );
  INVX1_RVT U14 ( .A(n70), .Y(n69) );
  INVX1_RVT U15 ( .A(\ab[10][23] ), .Y(n70) );
  INVX1_RVT U16 ( .A(n60), .Y(n59) );
  INVX1_RVT U17 ( .A(n66), .Y(n65) );
  INVX1_RVT U18 ( .A(\ab[8][23] ), .Y(n66) );
  INVX1_RVT U19 ( .A(n68), .Y(n67) );
  INVX1_RVT U20 ( .A(\ab[9][23] ), .Y(n68) );
  INVX1_RVT U21 ( .A(n56), .Y(n55) );
  INVX1_RVT U22 ( .A(\ab[3][23] ), .Y(n56) );
  INVX1_RVT U23 ( .A(n76), .Y(n75) );
  INVX1_RVT U24 ( .A(n64), .Y(n63) );
  INVX1_RVT U25 ( .A(\ab[7][23] ), .Y(n64) );
  INVX1_RVT U26 ( .A(n62), .Y(n61) );
  INVX1_RVT U27 ( .A(\ab[6][23] ), .Y(n62) );
  INVX1_RVT U28 ( .A(n54), .Y(n53) );
  INVX1_RVT U29 ( .A(\ab[2][23] ), .Y(n54) );
  INVX1_RVT U30 ( .A(n52), .Y(n51) );
  INVX1_RVT U31 ( .A(\ab[1][23] ), .Y(n52) );
  INVX1_RVT U32 ( .A(n50), .Y(n49) );
  INVX1_RVT U33 ( .A(\ab[0][23] ), .Y(n50) );
  XOR2X1_RVT U34 ( .A1(\CARRYB[23][11] ), .A2(\SUMB[23][12] ), .Y(\A1[33] ) );
  XOR2X1_RVT U35 ( .A1(\CARRYB[23][15] ), .A2(\SUMB[23][16] ), .Y(\A1[37] ) );
  XOR2X1_RVT U36 ( .A1(\CARRYB[23][5] ), .A2(\SUMB[23][6] ), .Y(\A1[27] ) );
  XOR2X1_RVT U37 ( .A1(\CARRYB[23][10] ), .A2(\SUMB[23][11] ), .Y(\A1[32] ) );
  XOR2X1_RVT U38 ( .A1(\CARRYB[23][9] ), .A2(\SUMB[23][10] ), .Y(\A1[31] ) );
  XOR2X1_RVT U39 ( .A1(\CARRYB[23][13] ), .A2(\SUMB[23][14] ), .Y(\A1[35] ) );
  XOR2X1_RVT U40 ( .A1(\CARRYB[23][14] ), .A2(\SUMB[23][15] ), .Y(\A1[36] ) );
  XOR2X1_RVT U41 ( .A1(\CARRYB[23][3] ), .A2(\SUMB[23][4] ), .Y(\A1[25] ) );
  XOR2X1_RVT U42 ( .A1(\CARRYB[23][7] ), .A2(\SUMB[23][8] ), .Y(\A1[29] ) );
  XOR2X1_RVT U43 ( .A1(\CARRYB[23][8] ), .A2(\SUMB[23][9] ), .Y(\A1[30] ) );
  XOR2X1_RVT U44 ( .A1(\CARRYB[23][4] ), .A2(\SUMB[23][5] ), .Y(\A1[26] ) );
  XOR2X1_RVT U45 ( .A1(\CARRYB[23][12] ), .A2(\SUMB[23][13] ), .Y(\A1[34] ) );
  XOR2X1_RVT U46 ( .A1(\CARRYB[23][6] ), .A2(\SUMB[23][7] ), .Y(\A1[28] ) );
  AND2X1_RVT U47 ( .A1(\CARRYB[23][11] ), .A2(\SUMB[23][12] ), .Y(\A2[34] ) );
  AND2X1_RVT U48 ( .A1(\CARRYB[23][15] ), .A2(\SUMB[23][16] ), .Y(\A2[38] ) );
  AND2X1_RVT U49 ( .A1(\CARRYB[23][5] ), .A2(\SUMB[23][6] ), .Y(\A2[28] ) );
  AND2X1_RVT U50 ( .A1(\CARRYB[23][10] ), .A2(\SUMB[23][11] ), .Y(\A2[33] ) );
  AND2X1_RVT U51 ( .A1(\CARRYB[23][9] ), .A2(\SUMB[23][10] ), .Y(\A2[32] ) );
  AND2X1_RVT U52 ( .A1(\CARRYB[23][13] ), .A2(\SUMB[23][14] ), .Y(\A2[36] ) );
  AND2X1_RVT U53 ( .A1(\CARRYB[23][14] ), .A2(\SUMB[23][15] ), .Y(\A2[37] ) );
  AND2X1_RVT U54 ( .A1(\CARRYB[23][7] ), .A2(\SUMB[23][8] ), .Y(\A2[30] ) );
  AND2X1_RVT U55 ( .A1(\CARRYB[23][3] ), .A2(\SUMB[23][4] ), .Y(\A2[26] ) );
  AND2X1_RVT U56 ( .A1(\CARRYB[23][8] ), .A2(\SUMB[23][9] ), .Y(\A2[31] ) );
  AND2X1_RVT U57 ( .A1(\CARRYB[23][4] ), .A2(\SUMB[23][5] ), .Y(\A2[27] ) );
  AND2X1_RVT U58 ( .A1(\CARRYB[23][12] ), .A2(\SUMB[23][13] ), .Y(\A2[35] ) );
  AND2X1_RVT U59 ( .A1(\CARRYB[23][6] ), .A2(\SUMB[23][7] ), .Y(\A2[29] ) );
  XOR2X1_RVT U60 ( .A1(\CARRYB[23][2] ), .A2(\SUMB[23][3] ), .Y(\A1[24] ) );
  AND2X1_RVT U61 ( .A1(\CARRYB[23][2] ), .A2(\SUMB[23][3] ), .Y(\A2[25] ) );
  XOR2X1_RVT U62 ( .A1(\CARRYB[23][1] ), .A2(\SUMB[23][2] ), .Y(\A1[23] ) );
  AND2X1_RVT U63 ( .A1(\CARRYB[23][1] ), .A2(\SUMB[23][2] ), .Y(\A2[24] ) );
  AND2X1_RVT U64 ( .A1(\CARRYB[23][0] ), .A2(\SUMB[23][1] ), .Y(\A2[23] ) );
  INVX1_RVT U65 ( .A(n90), .Y(n89) );
  INVX1_RVT U66 ( .A(n84), .Y(n83) );
  INVX1_RVT U67 ( .A(n88), .Y(n87) );
  INVX1_RVT U68 ( .A(\ab[19][23] ), .Y(n88) );
  INVX1_RVT U69 ( .A(n80), .Y(n79) );
  INVX1_RVT U70 ( .A(n86), .Y(n85) );
  INVX1_RVT U71 ( .A(n78), .Y(n77) );
  INVX1_RVT U72 ( .A(\ab[14][23] ), .Y(n78) );
  INVX1_RVT U73 ( .A(n82), .Y(n81) );
  XOR2X1_RVT U74 ( .A1(\CARRYB[23][19] ), .A2(\SUMB[23][20] ), .Y(\A1[41] ) );
  XOR2X1_RVT U75 ( .A1(\CARRYB[23][21] ), .A2(\SUMB[23][22] ), .Y(\A1[43] ) );
  XOR2X1_RVT U76 ( .A1(\CARRYB[23][18] ), .A2(\SUMB[23][19] ), .Y(\A1[40] ) );
  XOR2X1_RVT U77 ( .A1(\CARRYB[23][17] ), .A2(\SUMB[23][18] ), .Y(\A1[39] ) );
  XOR2X1_RVT U78 ( .A1(\CARRYB[23][20] ), .A2(\SUMB[23][21] ), .Y(\A1[42] ) );
  XOR2X1_RVT U79 ( .A1(\CARRYB[23][16] ), .A2(\SUMB[23][17] ), .Y(\A1[38] ) );
  AND2X1_RVT U80 ( .A1(\CARRYB[23][21] ), .A2(\SUMB[23][22] ), .Y(\A2[44] ) );
  AND2X1_RVT U81 ( .A1(\CARRYB[23][19] ), .A2(\SUMB[23][20] ), .Y(\A2[42] ) );
  AND2X1_RVT U82 ( .A1(\CARRYB[23][18] ), .A2(\SUMB[23][19] ), .Y(\A2[41] ) );
  AND2X1_RVT U83 ( .A1(\CARRYB[23][17] ), .A2(\SUMB[23][18] ), .Y(\A2[40] ) );
  AND2X1_RVT U84 ( .A1(\CARRYB[23][20] ), .A2(\SUMB[23][21] ), .Y(\A2[43] ) );
  AND2X1_RVT U85 ( .A1(\CARRYB[23][16] ), .A2(\SUMB[23][17] ), .Y(\A2[39] ) );
  INVX1_RVT U86 ( .A(n92), .Y(n91) );
  INVX1_RVT U87 ( .A(n94), .Y(n93) );
  INVX1_RVT U88 ( .A(\ab[22][23] ), .Y(n94) );
  INVX1_RVT U89 ( .A(\CARRYB[23][22] ), .Y(n95) );
  AND2X1_RVT U90 ( .A1(\ab[1][22] ), .A2(n49), .Y(\CARRYB[1][22] ) );
  AND2X1_RVT U91 ( .A1(\ab[1][21] ), .A2(\ab[0][22] ), .Y(\CARRYB[1][21] ) );
  XOR2X1_RVT U92 ( .A1(n49), .A2(\ab[1][22] ), .Y(\SUMB[1][22] ) );
  AND2X1_RVT U93 ( .A1(\ab[1][10] ), .A2(\ab[0][11] ), .Y(\CARRYB[1][10] ) );
  XOR2X1_RVT U94 ( .A1(\ab[0][12] ), .A2(\ab[1][11] ), .Y(\SUMB[1][11] ) );
  AND2X1_RVT U95 ( .A1(\ab[1][14] ), .A2(\ab[0][15] ), .Y(\CARRYB[1][14] ) );
  XOR2X1_RVT U96 ( .A1(\ab[0][16] ), .A2(\ab[1][15] ), .Y(\SUMB[1][15] ) );
  AND2X1_RVT U97 ( .A1(\ab[1][8] ), .A2(\ab[0][9] ), .Y(\CARRYB[1][8] ) );
  XOR2X1_RVT U98 ( .A1(\ab[0][10] ), .A2(\ab[1][9] ), .Y(\SUMB[1][9] ) );
  AND2X1_RVT U99 ( .A1(\ab[1][4] ), .A2(\ab[0][5] ), .Y(\CARRYB[1][4] ) );
  XOR2X1_RVT U100 ( .A1(\ab[0][6] ), .A2(\ab[1][5] ), .Y(\SUMB[1][5] ) );
  AND2X1_RVT U101 ( .A1(\ab[1][2] ), .A2(\ab[0][3] ), .Y(\CARRYB[1][2] ) );
  XOR2X1_RVT U102 ( .A1(\ab[0][4] ), .A2(\ab[1][3] ), .Y(\SUMB[1][3] ) );
  AND2X1_RVT U103 ( .A1(\ab[1][19] ), .A2(\ab[0][20] ), .Y(\CARRYB[1][19] ) );
  XOR2X1_RVT U104 ( .A1(\ab[0][21] ), .A2(\ab[1][20] ), .Y(\SUMB[1][20] ) );
  AND2X1_RVT U105 ( .A1(\ab[1][15] ), .A2(\ab[0][16] ), .Y(\CARRYB[1][15] ) );
  XOR2X1_RVT U106 ( .A1(\ab[0][17] ), .A2(\ab[1][16] ), .Y(\SUMB[1][16] ) );
  AND2X1_RVT U107 ( .A1(\ab[1][11] ), .A2(\ab[0][12] ), .Y(\CARRYB[1][11] ) );
  XOR2X1_RVT U108 ( .A1(\ab[0][13] ), .A2(\ab[1][12] ), .Y(\SUMB[1][12] ) );
  AND2X1_RVT U109 ( .A1(\ab[1][5] ), .A2(\ab[0][6] ), .Y(\CARRYB[1][5] ) );
  XOR2X1_RVT U110 ( .A1(\ab[0][7] ), .A2(\ab[1][6] ), .Y(\SUMB[1][6] ) );
  AND2X1_RVT U111 ( .A1(\ab[1][9] ), .A2(\ab[0][10] ), .Y(\CARRYB[1][9] ) );
  XOR2X1_RVT U112 ( .A1(\ab[0][11] ), .A2(\ab[1][10] ), .Y(\SUMB[1][10] ) );
  AND2X1_RVT U113 ( .A1(\ab[1][13] ), .A2(\ab[0][14] ), .Y(\CARRYB[1][13] ) );
  XOR2X1_RVT U114 ( .A1(\ab[0][15] ), .A2(\ab[1][14] ), .Y(\SUMB[1][14] ) );
  AND2X1_RVT U115 ( .A1(\ab[1][7] ), .A2(\ab[0][8] ), .Y(\CARRYB[1][7] ) );
  XOR2X1_RVT U116 ( .A1(\ab[0][9] ), .A2(\ab[1][8] ), .Y(\SUMB[1][8] ) );
  AND2X1_RVT U117 ( .A1(\ab[1][3] ), .A2(\ab[0][4] ), .Y(\CARRYB[1][3] ) );
  XOR2X1_RVT U118 ( .A1(\ab[0][5] ), .A2(\ab[1][4] ), .Y(\SUMB[1][4] ) );
  AND2X1_RVT U119 ( .A1(\ab[1][17] ), .A2(\ab[0][18] ), .Y(\CARRYB[1][17] ) );
  XOR2X1_RVT U120 ( .A1(\ab[0][19] ), .A2(\ab[1][18] ), .Y(\SUMB[1][18] ) );
  AND2X1_RVT U121 ( .A1(\ab[1][20] ), .A2(\ab[0][21] ), .Y(\CARRYB[1][20] ) );
  XOR2X1_RVT U122 ( .A1(\ab[0][22] ), .A2(\ab[1][21] ), .Y(\SUMB[1][21] ) );
  AND2X1_RVT U123 ( .A1(\ab[1][12] ), .A2(\ab[0][13] ), .Y(\CARRYB[1][12] ) );
  XOR2X1_RVT U124 ( .A1(\ab[0][14] ), .A2(\ab[1][13] ), .Y(\SUMB[1][13] ) );
  AND2X1_RVT U125 ( .A1(\ab[1][16] ), .A2(\ab[0][17] ), .Y(\CARRYB[1][16] ) );
  XOR2X1_RVT U126 ( .A1(\ab[0][18] ), .A2(\ab[1][17] ), .Y(\SUMB[1][17] ) );
  AND2X1_RVT U127 ( .A1(\ab[1][6] ), .A2(\ab[0][7] ), .Y(\CARRYB[1][6] ) );
  XOR2X1_RVT U128 ( .A1(\ab[0][8] ), .A2(\ab[1][7] ), .Y(\SUMB[1][7] ) );
  AND2X1_RVT U129 ( .A1(\ab[1][18] ), .A2(\ab[0][19] ), .Y(\CARRYB[1][18] ) );
  XOR2X1_RVT U130 ( .A1(\ab[0][20] ), .A2(\ab[1][19] ), .Y(\SUMB[1][19] ) );
  AND2X1_RVT U131 ( .A1(\ab[1][0] ), .A2(\ab[0][1] ), .Y(\CARRYB[1][0] ) );
  XOR2X1_RVT U132 ( .A1(\ab[0][2] ), .A2(\ab[1][1] ), .Y(\SUMB[1][1] ) );
  AND2X1_RVT U133 ( .A1(\ab[1][1] ), .A2(\ab[0][2] ), .Y(\CARRYB[1][1] ) );
  XOR2X1_RVT U134 ( .A1(\ab[0][3] ), .A2(\ab[1][2] ), .Y(\SUMB[1][2] ) );
  XOR2X1_RVT U135 ( .A1(\CARRYB[23][0] ), .A2(\SUMB[23][1] ), .Y(\A1[22] ) );
  XOR2X1_RVT U136 ( .A1(\ab[0][1] ), .A2(\ab[1][0] ), .Y(PRODUCT[1]) );
  INVX1_RVT U137 ( .A(n14), .Y(n13) );
  INVX1_RVT U138 ( .A(\ab[23][5] ), .Y(n14) );
  INVX1_RVT U139 ( .A(n42), .Y(n41) );
  INVX1_RVT U140 ( .A(\ab[23][19] ), .Y(n42) );
  INVX1_RVT U141 ( .A(n34), .Y(n33) );
  INVX1_RVT U142 ( .A(\ab[23][15] ), .Y(n34) );
  INVX1_RVT U143 ( .A(n26), .Y(n25) );
  INVX1_RVT U144 ( .A(\ab[23][11] ), .Y(n26) );
  INVX1_RVT U145 ( .A(n46), .Y(n45) );
  INVX1_RVT U146 ( .A(\ab[23][21] ), .Y(n46) );
  INVX1_RVT U147 ( .A(n24), .Y(n23) );
  INVX1_RVT U148 ( .A(\ab[23][10] ), .Y(n24) );
  INVX1_RVT U149 ( .A(n40), .Y(n39) );
  INVX1_RVT U150 ( .A(\ab[23][18] ), .Y(n40) );
  INVX1_RVT U151 ( .A(n48), .Y(n47) );
  INVX1_RVT U152 ( .A(\ab[23][22] ), .Y(n48) );
  INVX1_RVT U153 ( .A(n22), .Y(n21) );
  INVX1_RVT U154 ( .A(\ab[23][9] ), .Y(n22) );
  INVX1_RVT U155 ( .A(n30), .Y(n29) );
  INVX1_RVT U156 ( .A(\ab[23][13] ), .Y(n30) );
  INVX1_RVT U157 ( .A(n32), .Y(n31) );
  INVX1_RVT U158 ( .A(\ab[23][14] ), .Y(n32) );
  INVX1_RVT U159 ( .A(n38), .Y(n37) );
  INVX1_RVT U160 ( .A(\ab[23][17] ), .Y(n38) );
  INVX1_RVT U161 ( .A(n18), .Y(n17) );
  INVX1_RVT U162 ( .A(\ab[23][7] ), .Y(n18) );
  INVX1_RVT U163 ( .A(n10), .Y(n9) );
  INVX1_RVT U164 ( .A(\ab[23][3] ), .Y(n10) );
  INVX1_RVT U165 ( .A(n20), .Y(n19) );
  INVX1_RVT U166 ( .A(\ab[23][8] ), .Y(n20) );
  INVX1_RVT U167 ( .A(n12), .Y(n11) );
  INVX1_RVT U168 ( .A(\ab[23][4] ), .Y(n12) );
  INVX1_RVT U169 ( .A(n44), .Y(n43) );
  INVX1_RVT U170 ( .A(\ab[23][20] ), .Y(n44) );
  INVX1_RVT U171 ( .A(n28), .Y(n27) );
  INVX1_RVT U172 ( .A(\ab[23][12] ), .Y(n28) );
  INVX1_RVT U173 ( .A(n36), .Y(n35) );
  INVX1_RVT U174 ( .A(\ab[23][16] ), .Y(n36) );
  INVX1_RVT U175 ( .A(n16), .Y(n15) );
  INVX1_RVT U176 ( .A(\ab[23][6] ), .Y(n16) );
  INVX1_RVT U177 ( .A(n72), .Y(n71) );
  INVX1_RVT U178 ( .A(n8), .Y(n7) );
  INVX1_RVT U179 ( .A(\ab[23][2] ), .Y(n8) );
  INVX1_RVT U180 ( .A(n6), .Y(n5) );
  INVX1_RVT U181 ( .A(\ab[23][1] ), .Y(n6) );
  INVX1_RVT U182 ( .A(n4), .Y(n3) );
  INVX1_RVT U183 ( .A(\ab[23][0] ), .Y(n4) );
  INVX0_RVT U184 ( .A(\ab[21][23] ), .Y(n92) );
  AND2X1_RVT U186 ( .A1(n21), .A2(n67), .Y(\ab[9][9] ) );
  AND2X1_RVT U187 ( .A1(n19), .A2(n67), .Y(\ab[9][8] ) );
  AND2X1_RVT U188 ( .A1(n17), .A2(n67), .Y(\ab[9][7] ) );
  AND2X1_RVT U189 ( .A1(n15), .A2(n67), .Y(\ab[9][6] ) );
  AND2X1_RVT U190 ( .A1(n13), .A2(n67), .Y(\ab[9][5] ) );
  AND2X1_RVT U191 ( .A1(n11), .A2(n67), .Y(\ab[9][4] ) );
  AND2X1_RVT U192 ( .A1(n9), .A2(n67), .Y(\ab[9][3] ) );
  AND2X1_RVT U193 ( .A1(n7), .A2(n67), .Y(\ab[9][2] ) );
  AND2X1_RVT U194 ( .A1(n47), .A2(n67), .Y(\ab[9][22] ) );
  AND2X1_RVT U195 ( .A1(n45), .A2(n67), .Y(\ab[9][21] ) );
  AND2X1_RVT U196 ( .A1(n43), .A2(n67), .Y(\ab[9][20] ) );
  AND2X1_RVT U197 ( .A1(n5), .A2(n67), .Y(\ab[9][1] ) );
  AND2X1_RVT U198 ( .A1(n41), .A2(n67), .Y(\ab[9][19] ) );
  AND2X1_RVT U199 ( .A1(n39), .A2(n67), .Y(\ab[9][18] ) );
  AND2X1_RVT U200 ( .A1(n37), .A2(n67), .Y(\ab[9][17] ) );
  AND2X1_RVT U201 ( .A1(n35), .A2(n67), .Y(\ab[9][16] ) );
  AND2X1_RVT U202 ( .A1(n33), .A2(n67), .Y(\ab[9][15] ) );
  AND2X1_RVT U203 ( .A1(n31), .A2(n67), .Y(\ab[9][14] ) );
  AND2X1_RVT U204 ( .A1(n29), .A2(n67), .Y(\ab[9][13] ) );
  AND2X1_RVT U205 ( .A1(n27), .A2(n67), .Y(\ab[9][12] ) );
  AND2X1_RVT U206 ( .A1(n25), .A2(n67), .Y(\ab[9][11] ) );
  AND2X1_RVT U207 ( .A1(n23), .A2(n67), .Y(\ab[9][10] ) );
  AND2X1_RVT U208 ( .A1(n3), .A2(n67), .Y(\ab[9][0] ) );
  AND2X1_RVT U209 ( .A1(n65), .A2(n21), .Y(\ab[8][9] ) );
  AND2X1_RVT U210 ( .A1(n65), .A2(n19), .Y(\ab[8][8] ) );
  AND2X1_RVT U211 ( .A1(n65), .A2(n17), .Y(\ab[8][7] ) );
  AND2X1_RVT U212 ( .A1(n65), .A2(n15), .Y(\ab[8][6] ) );
  AND2X1_RVT U213 ( .A1(n65), .A2(n13), .Y(\ab[8][5] ) );
  AND2X1_RVT U214 ( .A1(n65), .A2(n11), .Y(\ab[8][4] ) );
  AND2X1_RVT U215 ( .A1(n65), .A2(n9), .Y(\ab[8][3] ) );
  AND2X1_RVT U216 ( .A1(n65), .A2(n7), .Y(\ab[8][2] ) );
  AND2X1_RVT U217 ( .A1(n65), .A2(n47), .Y(\ab[8][22] ) );
  AND2X1_RVT U218 ( .A1(n65), .A2(n45), .Y(\ab[8][21] ) );
  AND2X1_RVT U219 ( .A1(n65), .A2(n43), .Y(\ab[8][20] ) );
  AND2X1_RVT U220 ( .A1(n65), .A2(n5), .Y(\ab[8][1] ) );
  AND2X1_RVT U221 ( .A1(n65), .A2(n41), .Y(\ab[8][19] ) );
  AND2X1_RVT U222 ( .A1(n65), .A2(n39), .Y(\ab[8][18] ) );
  AND2X1_RVT U223 ( .A1(n65), .A2(n37), .Y(\ab[8][17] ) );
  AND2X1_RVT U224 ( .A1(n65), .A2(n35), .Y(\ab[8][16] ) );
  AND2X1_RVT U225 ( .A1(n65), .A2(n33), .Y(\ab[8][15] ) );
  AND2X1_RVT U226 ( .A1(n65), .A2(n31), .Y(\ab[8][14] ) );
  AND2X1_RVT U227 ( .A1(n65), .A2(n29), .Y(\ab[8][13] ) );
  AND2X1_RVT U228 ( .A1(n65), .A2(n27), .Y(\ab[8][12] ) );
  AND2X1_RVT U229 ( .A1(n65), .A2(n25), .Y(\ab[8][11] ) );
  AND2X1_RVT U230 ( .A1(n65), .A2(n23), .Y(\ab[8][10] ) );
  AND2X1_RVT U231 ( .A1(n65), .A2(n3), .Y(\ab[8][0] ) );
  AND2X1_RVT U232 ( .A1(n63), .A2(n21), .Y(\ab[7][9] ) );
  AND2X1_RVT U233 ( .A1(n63), .A2(n19), .Y(\ab[7][8] ) );
  AND2X1_RVT U234 ( .A1(n63), .A2(n17), .Y(\ab[7][7] ) );
  AND2X1_RVT U235 ( .A1(n63), .A2(n15), .Y(\ab[7][6] ) );
  AND2X1_RVT U236 ( .A1(n63), .A2(n13), .Y(\ab[7][5] ) );
  AND2X1_RVT U237 ( .A1(n63), .A2(n11), .Y(\ab[7][4] ) );
  AND2X1_RVT U238 ( .A1(n63), .A2(n9), .Y(\ab[7][3] ) );
  AND2X1_RVT U239 ( .A1(n63), .A2(n7), .Y(\ab[7][2] ) );
  AND2X1_RVT U240 ( .A1(n63), .A2(n47), .Y(\ab[7][22] ) );
  AND2X1_RVT U241 ( .A1(n63), .A2(n45), .Y(\ab[7][21] ) );
  AND2X1_RVT U242 ( .A1(n63), .A2(n43), .Y(\ab[7][20] ) );
  AND2X1_RVT U243 ( .A1(n63), .A2(n5), .Y(\ab[7][1] ) );
  AND2X1_RVT U244 ( .A1(n63), .A2(n41), .Y(\ab[7][19] ) );
  AND2X1_RVT U245 ( .A1(n63), .A2(n39), .Y(\ab[7][18] ) );
  AND2X1_RVT U246 ( .A1(n63), .A2(n37), .Y(\ab[7][17] ) );
  AND2X1_RVT U247 ( .A1(n63), .A2(n35), .Y(\ab[7][16] ) );
  AND2X1_RVT U248 ( .A1(n63), .A2(n33), .Y(\ab[7][15] ) );
  AND2X1_RVT U249 ( .A1(n63), .A2(n31), .Y(\ab[7][14] ) );
  AND2X1_RVT U250 ( .A1(n63), .A2(n29), .Y(\ab[7][13] ) );
  AND2X1_RVT U251 ( .A1(n63), .A2(n27), .Y(\ab[7][12] ) );
  AND2X1_RVT U252 ( .A1(n63), .A2(n25), .Y(\ab[7][11] ) );
  AND2X1_RVT U253 ( .A1(n63), .A2(n23), .Y(\ab[7][10] ) );
  AND2X1_RVT U254 ( .A1(n63), .A2(n3), .Y(\ab[7][0] ) );
  AND2X1_RVT U255 ( .A1(n61), .A2(n21), .Y(\ab[6][9] ) );
  AND2X1_RVT U256 ( .A1(n61), .A2(n19), .Y(\ab[6][8] ) );
  AND2X1_RVT U257 ( .A1(n61), .A2(n17), .Y(\ab[6][7] ) );
  AND2X1_RVT U258 ( .A1(n61), .A2(n15), .Y(\ab[6][6] ) );
  AND2X1_RVT U259 ( .A1(n61), .A2(n13), .Y(\ab[6][5] ) );
  AND2X1_RVT U260 ( .A1(n61), .A2(n11), .Y(\ab[6][4] ) );
  AND2X1_RVT U261 ( .A1(n61), .A2(n9), .Y(\ab[6][3] ) );
  AND2X1_RVT U262 ( .A1(n61), .A2(n7), .Y(\ab[6][2] ) );
  AND2X1_RVT U263 ( .A1(n61), .A2(n47), .Y(\ab[6][22] ) );
  AND2X1_RVT U264 ( .A1(n61), .A2(n45), .Y(\ab[6][21] ) );
  AND2X1_RVT U265 ( .A1(n61), .A2(n43), .Y(\ab[6][20] ) );
  AND2X1_RVT U266 ( .A1(n61), .A2(n5), .Y(\ab[6][1] ) );
  AND2X1_RVT U267 ( .A1(n61), .A2(n41), .Y(\ab[6][19] ) );
  AND2X1_RVT U268 ( .A1(n61), .A2(n39), .Y(\ab[6][18] ) );
  AND2X1_RVT U269 ( .A1(n61), .A2(n37), .Y(\ab[6][17] ) );
  AND2X1_RVT U270 ( .A1(n61), .A2(n35), .Y(\ab[6][16] ) );
  AND2X1_RVT U271 ( .A1(n61), .A2(n33), .Y(\ab[6][15] ) );
  AND2X1_RVT U272 ( .A1(n61), .A2(n31), .Y(\ab[6][14] ) );
  AND2X1_RVT U273 ( .A1(n61), .A2(n29), .Y(\ab[6][13] ) );
  AND2X1_RVT U274 ( .A1(n61), .A2(n27), .Y(\ab[6][12] ) );
  AND2X1_RVT U275 ( .A1(n61), .A2(n25), .Y(\ab[6][11] ) );
  AND2X1_RVT U276 ( .A1(n61), .A2(n23), .Y(\ab[6][10] ) );
  AND2X1_RVT U277 ( .A1(n61), .A2(n3), .Y(\ab[6][0] ) );
  AND2X1_RVT U278 ( .A1(n59), .A2(n21), .Y(\ab[5][9] ) );
  AND2X1_RVT U279 ( .A1(n59), .A2(n19), .Y(\ab[5][8] ) );
  AND2X1_RVT U280 ( .A1(n59), .A2(n17), .Y(\ab[5][7] ) );
  AND2X1_RVT U281 ( .A1(n59), .A2(n15), .Y(\ab[5][6] ) );
  AND2X1_RVT U282 ( .A1(n59), .A2(n13), .Y(\ab[5][5] ) );
  AND2X1_RVT U283 ( .A1(n59), .A2(n11), .Y(\ab[5][4] ) );
  AND2X1_RVT U284 ( .A1(n59), .A2(n9), .Y(\ab[5][3] ) );
  AND2X1_RVT U285 ( .A1(n59), .A2(n7), .Y(\ab[5][2] ) );
  AND2X1_RVT U286 ( .A1(n59), .A2(n47), .Y(\ab[5][22] ) );
  AND2X1_RVT U287 ( .A1(n59), .A2(n45), .Y(\ab[5][21] ) );
  AND2X1_RVT U288 ( .A1(n59), .A2(n43), .Y(\ab[5][20] ) );
  AND2X1_RVT U289 ( .A1(n59), .A2(n5), .Y(\ab[5][1] ) );
  AND2X1_RVT U290 ( .A1(n59), .A2(n41), .Y(\ab[5][19] ) );
  AND2X1_RVT U291 ( .A1(n59), .A2(n39), .Y(\ab[5][18] ) );
  AND2X1_RVT U292 ( .A1(n59), .A2(n37), .Y(\ab[5][17] ) );
  AND2X1_RVT U293 ( .A1(n59), .A2(n35), .Y(\ab[5][16] ) );
  AND2X1_RVT U294 ( .A1(n59), .A2(n33), .Y(\ab[5][15] ) );
  AND2X1_RVT U295 ( .A1(n59), .A2(n31), .Y(\ab[5][14] ) );
  AND2X1_RVT U296 ( .A1(n59), .A2(n29), .Y(\ab[5][13] ) );
  AND2X1_RVT U297 ( .A1(n59), .A2(n27), .Y(\ab[5][12] ) );
  AND2X1_RVT U298 ( .A1(n59), .A2(n25), .Y(\ab[5][11] ) );
  AND2X1_RVT U299 ( .A1(n59), .A2(n23), .Y(\ab[5][10] ) );
  AND2X1_RVT U300 ( .A1(n59), .A2(n3), .Y(\ab[5][0] ) );
  AND2X1_RVT U301 ( .A1(n57), .A2(n21), .Y(\ab[4][9] ) );
  AND2X1_RVT U302 ( .A1(n57), .A2(n19), .Y(\ab[4][8] ) );
  AND2X1_RVT U303 ( .A1(n57), .A2(n17), .Y(\ab[4][7] ) );
  AND2X1_RVT U304 ( .A1(n57), .A2(n15), .Y(\ab[4][6] ) );
  AND2X1_RVT U305 ( .A1(n57), .A2(n13), .Y(\ab[4][5] ) );
  AND2X1_RVT U306 ( .A1(n57), .A2(n11), .Y(\ab[4][4] ) );
  AND2X1_RVT U307 ( .A1(n57), .A2(n9), .Y(\ab[4][3] ) );
  AND2X1_RVT U308 ( .A1(n57), .A2(n7), .Y(\ab[4][2] ) );
  AND2X1_RVT U309 ( .A1(n57), .A2(n47), .Y(\ab[4][22] ) );
  AND2X1_RVT U310 ( .A1(n57), .A2(n45), .Y(\ab[4][21] ) );
  AND2X1_RVT U311 ( .A1(n57), .A2(n43), .Y(\ab[4][20] ) );
  AND2X1_RVT U312 ( .A1(n57), .A2(n5), .Y(\ab[4][1] ) );
  AND2X1_RVT U313 ( .A1(n57), .A2(n41), .Y(\ab[4][19] ) );
  AND2X1_RVT U314 ( .A1(n57), .A2(n39), .Y(\ab[4][18] ) );
  AND2X1_RVT U315 ( .A1(n57), .A2(n37), .Y(\ab[4][17] ) );
  AND2X1_RVT U316 ( .A1(n57), .A2(n35), .Y(\ab[4][16] ) );
  AND2X1_RVT U317 ( .A1(n57), .A2(n33), .Y(\ab[4][15] ) );
  AND2X1_RVT U318 ( .A1(n57), .A2(n31), .Y(\ab[4][14] ) );
  AND2X1_RVT U319 ( .A1(n57), .A2(n29), .Y(\ab[4][13] ) );
  AND2X1_RVT U320 ( .A1(n57), .A2(n27), .Y(\ab[4][12] ) );
  AND2X1_RVT U321 ( .A1(n57), .A2(n25), .Y(\ab[4][11] ) );
  AND2X1_RVT U322 ( .A1(n57), .A2(n23), .Y(\ab[4][10] ) );
  AND2X1_RVT U323 ( .A1(n57), .A2(n3), .Y(\ab[4][0] ) );
  AND2X1_RVT U324 ( .A1(n55), .A2(n21), .Y(\ab[3][9] ) );
  AND2X1_RVT U325 ( .A1(n55), .A2(n19), .Y(\ab[3][8] ) );
  AND2X1_RVT U326 ( .A1(n55), .A2(n17), .Y(\ab[3][7] ) );
  AND2X1_RVT U327 ( .A1(n55), .A2(n15), .Y(\ab[3][6] ) );
  AND2X1_RVT U328 ( .A1(n55), .A2(n13), .Y(\ab[3][5] ) );
  AND2X1_RVT U329 ( .A1(n55), .A2(n11), .Y(\ab[3][4] ) );
  AND2X1_RVT U330 ( .A1(n55), .A2(n9), .Y(\ab[3][3] ) );
  AND2X1_RVT U331 ( .A1(n55), .A2(n7), .Y(\ab[3][2] ) );
  AND2X1_RVT U332 ( .A1(n55), .A2(n47), .Y(\ab[3][22] ) );
  AND2X1_RVT U333 ( .A1(n55), .A2(n45), .Y(\ab[3][21] ) );
  AND2X1_RVT U334 ( .A1(n55), .A2(n43), .Y(\ab[3][20] ) );
  AND2X1_RVT U335 ( .A1(n55), .A2(n5), .Y(\ab[3][1] ) );
  AND2X1_RVT U336 ( .A1(n55), .A2(n41), .Y(\ab[3][19] ) );
  AND2X1_RVT U337 ( .A1(n55), .A2(n39), .Y(\ab[3][18] ) );
  AND2X1_RVT U338 ( .A1(n55), .A2(n37), .Y(\ab[3][17] ) );
  AND2X1_RVT U339 ( .A1(n55), .A2(n35), .Y(\ab[3][16] ) );
  AND2X1_RVT U340 ( .A1(n55), .A2(n33), .Y(\ab[3][15] ) );
  AND2X1_RVT U341 ( .A1(n55), .A2(n31), .Y(\ab[3][14] ) );
  AND2X1_RVT U342 ( .A1(n55), .A2(n29), .Y(\ab[3][13] ) );
  AND2X1_RVT U343 ( .A1(n55), .A2(n27), .Y(\ab[3][12] ) );
  AND2X1_RVT U344 ( .A1(n55), .A2(n25), .Y(\ab[3][11] ) );
  AND2X1_RVT U345 ( .A1(n55), .A2(n23), .Y(\ab[3][10] ) );
  AND2X1_RVT U346 ( .A1(n55), .A2(n3), .Y(\ab[3][0] ) );
  AND2X1_RVT U347 ( .A1(n53), .A2(n21), .Y(\ab[2][9] ) );
  AND2X1_RVT U348 ( .A1(n53), .A2(n19), .Y(\ab[2][8] ) );
  AND2X1_RVT U349 ( .A1(n53), .A2(n17), .Y(\ab[2][7] ) );
  AND2X1_RVT U350 ( .A1(n53), .A2(n15), .Y(\ab[2][6] ) );
  AND2X1_RVT U351 ( .A1(n53), .A2(n13), .Y(\ab[2][5] ) );
  AND2X1_RVT U352 ( .A1(n53), .A2(n11), .Y(\ab[2][4] ) );
  AND2X1_RVT U353 ( .A1(n53), .A2(n9), .Y(\ab[2][3] ) );
  AND2X1_RVT U354 ( .A1(n53), .A2(n7), .Y(\ab[2][2] ) );
  AND2X1_RVT U355 ( .A1(n53), .A2(n47), .Y(\ab[2][22] ) );
  AND2X1_RVT U356 ( .A1(n53), .A2(n45), .Y(\ab[2][21] ) );
  AND2X1_RVT U357 ( .A1(n53), .A2(n43), .Y(\ab[2][20] ) );
  AND2X1_RVT U358 ( .A1(n53), .A2(n5), .Y(\ab[2][1] ) );
  AND2X1_RVT U359 ( .A1(n53), .A2(n41), .Y(\ab[2][19] ) );
  AND2X1_RVT U360 ( .A1(n53), .A2(n39), .Y(\ab[2][18] ) );
  AND2X1_RVT U361 ( .A1(n53), .A2(n37), .Y(\ab[2][17] ) );
  AND2X1_RVT U362 ( .A1(n53), .A2(n35), .Y(\ab[2][16] ) );
  AND2X1_RVT U363 ( .A1(n53), .A2(n33), .Y(\ab[2][15] ) );
  AND2X1_RVT U364 ( .A1(n53), .A2(n31), .Y(\ab[2][14] ) );
  AND2X1_RVT U365 ( .A1(n53), .A2(n29), .Y(\ab[2][13] ) );
  AND2X1_RVT U366 ( .A1(n53), .A2(n27), .Y(\ab[2][12] ) );
  AND2X1_RVT U367 ( .A1(n53), .A2(n25), .Y(\ab[2][11] ) );
  AND2X1_RVT U368 ( .A1(n53), .A2(n23), .Y(\ab[2][10] ) );
  AND2X1_RVT U369 ( .A1(n53), .A2(n3), .Y(\ab[2][0] ) );
  AND2X1_RVT U370 ( .A1(n93), .A2(n21), .Y(\ab[22][9] ) );
  AND2X1_RVT U371 ( .A1(n93), .A2(n19), .Y(\ab[22][8] ) );
  AND2X1_RVT U372 ( .A1(n93), .A2(n17), .Y(\ab[22][7] ) );
  AND2X1_RVT U373 ( .A1(n93), .A2(n15), .Y(\ab[22][6] ) );
  AND2X1_RVT U374 ( .A1(n93), .A2(n13), .Y(\ab[22][5] ) );
  AND2X1_RVT U375 ( .A1(n93), .A2(n11), .Y(\ab[22][4] ) );
  AND2X1_RVT U376 ( .A1(n93), .A2(n9), .Y(\ab[22][3] ) );
  AND2X1_RVT U377 ( .A1(n93), .A2(n7), .Y(\ab[22][2] ) );
  AND2X1_RVT U378 ( .A1(n93), .A2(n47), .Y(\ab[22][22] ) );
  AND2X1_RVT U379 ( .A1(n93), .A2(n45), .Y(\ab[22][21] ) );
  AND2X1_RVT U380 ( .A1(n93), .A2(n43), .Y(\ab[22][20] ) );
  AND2X1_RVT U381 ( .A1(n93), .A2(n5), .Y(\ab[22][1] ) );
  AND2X1_RVT U382 ( .A1(n93), .A2(n41), .Y(\ab[22][19] ) );
  AND2X1_RVT U383 ( .A1(n93), .A2(n39), .Y(\ab[22][18] ) );
  AND2X1_RVT U384 ( .A1(n93), .A2(n37), .Y(\ab[22][17] ) );
  AND2X1_RVT U385 ( .A1(n93), .A2(n35), .Y(\ab[22][16] ) );
  AND2X1_RVT U386 ( .A1(n93), .A2(n33), .Y(\ab[22][15] ) );
  AND2X1_RVT U387 ( .A1(n93), .A2(n31), .Y(\ab[22][14] ) );
  AND2X1_RVT U388 ( .A1(n93), .A2(n29), .Y(\ab[22][13] ) );
  AND2X1_RVT U389 ( .A1(n93), .A2(n27), .Y(\ab[22][12] ) );
  AND2X1_RVT U390 ( .A1(n93), .A2(n25), .Y(\ab[22][11] ) );
  AND2X1_RVT U391 ( .A1(n93), .A2(n23), .Y(\ab[22][10] ) );
  AND2X1_RVT U392 ( .A1(n93), .A2(n3), .Y(\ab[22][0] ) );
  AND2X1_RVT U393 ( .A1(n91), .A2(n21), .Y(\ab[21][9] ) );
  AND2X1_RVT U394 ( .A1(n91), .A2(n19), .Y(\ab[21][8] ) );
  AND2X1_RVT U395 ( .A1(n91), .A2(n17), .Y(\ab[21][7] ) );
  AND2X1_RVT U396 ( .A1(n91), .A2(n15), .Y(\ab[21][6] ) );
  AND2X1_RVT U397 ( .A1(n91), .A2(n13), .Y(\ab[21][5] ) );
  AND2X1_RVT U398 ( .A1(n91), .A2(n11), .Y(\ab[21][4] ) );
  AND2X1_RVT U399 ( .A1(n91), .A2(n9), .Y(\ab[21][3] ) );
  AND2X1_RVT U400 ( .A1(n91), .A2(n7), .Y(\ab[21][2] ) );
  AND2X1_RVT U401 ( .A1(n91), .A2(n47), .Y(\ab[21][22] ) );
  AND2X1_RVT U402 ( .A1(n91), .A2(n45), .Y(\ab[21][21] ) );
  AND2X1_RVT U403 ( .A1(n91), .A2(n43), .Y(\ab[21][20] ) );
  AND2X1_RVT U404 ( .A1(n91), .A2(n5), .Y(\ab[21][1] ) );
  AND2X1_RVT U405 ( .A1(n91), .A2(n41), .Y(\ab[21][19] ) );
  AND2X1_RVT U406 ( .A1(n91), .A2(n39), .Y(\ab[21][18] ) );
  AND2X1_RVT U407 ( .A1(n91), .A2(n37), .Y(\ab[21][17] ) );
  AND2X1_RVT U408 ( .A1(n91), .A2(n35), .Y(\ab[21][16] ) );
  AND2X1_RVT U409 ( .A1(n91), .A2(n33), .Y(\ab[21][15] ) );
  AND2X1_RVT U410 ( .A1(n91), .A2(n31), .Y(\ab[21][14] ) );
  AND2X1_RVT U411 ( .A1(n91), .A2(n29), .Y(\ab[21][13] ) );
  AND2X1_RVT U412 ( .A1(n91), .A2(n27), .Y(\ab[21][12] ) );
  AND2X1_RVT U413 ( .A1(n91), .A2(n25), .Y(\ab[21][11] ) );
  AND2X1_RVT U414 ( .A1(n91), .A2(n23), .Y(\ab[21][10] ) );
  AND2X1_RVT U415 ( .A1(n91), .A2(n3), .Y(\ab[21][0] ) );
  AND2X1_RVT U416 ( .A1(n89), .A2(n21), .Y(\ab[20][9] ) );
  AND2X1_RVT U417 ( .A1(n89), .A2(n19), .Y(\ab[20][8] ) );
  AND2X1_RVT U418 ( .A1(n89), .A2(n17), .Y(\ab[20][7] ) );
  AND2X1_RVT U419 ( .A1(n89), .A2(n15), .Y(\ab[20][6] ) );
  AND2X1_RVT U420 ( .A1(n89), .A2(n13), .Y(\ab[20][5] ) );
  AND2X1_RVT U421 ( .A1(n89), .A2(n11), .Y(\ab[20][4] ) );
  AND2X1_RVT U422 ( .A1(n89), .A2(n9), .Y(\ab[20][3] ) );
  AND2X1_RVT U423 ( .A1(n89), .A2(n7), .Y(\ab[20][2] ) );
  AND2X1_RVT U424 ( .A1(n89), .A2(n47), .Y(\ab[20][22] ) );
  AND2X1_RVT U425 ( .A1(n89), .A2(n45), .Y(\ab[20][21] ) );
  AND2X1_RVT U426 ( .A1(n89), .A2(n43), .Y(\ab[20][20] ) );
  AND2X1_RVT U427 ( .A1(n89), .A2(n5), .Y(\ab[20][1] ) );
  AND2X1_RVT U428 ( .A1(n89), .A2(n41), .Y(\ab[20][19] ) );
  AND2X1_RVT U429 ( .A1(n89), .A2(n39), .Y(\ab[20][18] ) );
  AND2X1_RVT U430 ( .A1(n89), .A2(n37), .Y(\ab[20][17] ) );
  AND2X1_RVT U431 ( .A1(n89), .A2(n35), .Y(\ab[20][16] ) );
  AND2X1_RVT U432 ( .A1(n89), .A2(n33), .Y(\ab[20][15] ) );
  AND2X1_RVT U433 ( .A1(n89), .A2(n31), .Y(\ab[20][14] ) );
  AND2X1_RVT U434 ( .A1(n89), .A2(n29), .Y(\ab[20][13] ) );
  AND2X1_RVT U435 ( .A1(n89), .A2(n27), .Y(\ab[20][12] ) );
  AND2X1_RVT U436 ( .A1(n89), .A2(n25), .Y(\ab[20][11] ) );
  AND2X1_RVT U437 ( .A1(n89), .A2(n23), .Y(\ab[20][10] ) );
  AND2X1_RVT U438 ( .A1(n89), .A2(n3), .Y(\ab[20][0] ) );
  AND2X1_RVT U439 ( .A1(n51), .A2(n21), .Y(\ab[1][9] ) );
  AND2X1_RVT U440 ( .A1(n51), .A2(n19), .Y(\ab[1][8] ) );
  AND2X1_RVT U441 ( .A1(n51), .A2(n17), .Y(\ab[1][7] ) );
  AND2X1_RVT U442 ( .A1(n51), .A2(n15), .Y(\ab[1][6] ) );
  AND2X1_RVT U443 ( .A1(n51), .A2(n13), .Y(\ab[1][5] ) );
  AND2X1_RVT U444 ( .A1(n51), .A2(n11), .Y(\ab[1][4] ) );
  AND2X1_RVT U445 ( .A1(n51), .A2(n9), .Y(\ab[1][3] ) );
  AND2X1_RVT U446 ( .A1(n51), .A2(n7), .Y(\ab[1][2] ) );
  AND2X1_RVT U447 ( .A1(n51), .A2(n47), .Y(\ab[1][22] ) );
  AND2X1_RVT U448 ( .A1(n51), .A2(n45), .Y(\ab[1][21] ) );
  AND2X1_RVT U449 ( .A1(n51), .A2(n43), .Y(\ab[1][20] ) );
  AND2X1_RVT U450 ( .A1(n51), .A2(n5), .Y(\ab[1][1] ) );
  AND2X1_RVT U451 ( .A1(n51), .A2(n41), .Y(\ab[1][19] ) );
  AND2X1_RVT U452 ( .A1(n51), .A2(n39), .Y(\ab[1][18] ) );
  AND2X1_RVT U453 ( .A1(n51), .A2(n37), .Y(\ab[1][17] ) );
  AND2X1_RVT U454 ( .A1(n51), .A2(n35), .Y(\ab[1][16] ) );
  AND2X1_RVT U455 ( .A1(n51), .A2(n33), .Y(\ab[1][15] ) );
  AND2X1_RVT U456 ( .A1(n51), .A2(n31), .Y(\ab[1][14] ) );
  AND2X1_RVT U457 ( .A1(n51), .A2(n29), .Y(\ab[1][13] ) );
  AND2X1_RVT U458 ( .A1(n51), .A2(n27), .Y(\ab[1][12] ) );
  AND2X1_RVT U459 ( .A1(n51), .A2(n25), .Y(\ab[1][11] ) );
  AND2X1_RVT U460 ( .A1(n51), .A2(n23), .Y(\ab[1][10] ) );
  AND2X1_RVT U461 ( .A1(n51), .A2(n3), .Y(\ab[1][0] ) );
  AND2X1_RVT U462 ( .A1(n87), .A2(n21), .Y(\ab[19][9] ) );
  AND2X1_RVT U463 ( .A1(n87), .A2(n19), .Y(\ab[19][8] ) );
  AND2X1_RVT U464 ( .A1(n87), .A2(n17), .Y(\ab[19][7] ) );
  AND2X1_RVT U465 ( .A1(n87), .A2(n15), .Y(\ab[19][6] ) );
  AND2X1_RVT U466 ( .A1(n87), .A2(n13), .Y(\ab[19][5] ) );
  AND2X1_RVT U467 ( .A1(n87), .A2(n11), .Y(\ab[19][4] ) );
  AND2X1_RVT U468 ( .A1(n87), .A2(n9), .Y(\ab[19][3] ) );
  AND2X1_RVT U469 ( .A1(n87), .A2(n7), .Y(\ab[19][2] ) );
  AND2X1_RVT U470 ( .A1(n87), .A2(n47), .Y(\ab[19][22] ) );
  AND2X1_RVT U471 ( .A1(n87), .A2(n45), .Y(\ab[19][21] ) );
  AND2X1_RVT U472 ( .A1(n87), .A2(n43), .Y(\ab[19][20] ) );
  AND2X1_RVT U473 ( .A1(n87), .A2(n5), .Y(\ab[19][1] ) );
  AND2X1_RVT U474 ( .A1(n87), .A2(n41), .Y(\ab[19][19] ) );
  AND2X1_RVT U475 ( .A1(n87), .A2(n39), .Y(\ab[19][18] ) );
  AND2X1_RVT U476 ( .A1(n87), .A2(n37), .Y(\ab[19][17] ) );
  AND2X1_RVT U477 ( .A1(n87), .A2(n35), .Y(\ab[19][16] ) );
  AND2X1_RVT U478 ( .A1(n87), .A2(n33), .Y(\ab[19][15] ) );
  AND2X1_RVT U479 ( .A1(n87), .A2(n31), .Y(\ab[19][14] ) );
  AND2X1_RVT U480 ( .A1(n87), .A2(n29), .Y(\ab[19][13] ) );
  AND2X1_RVT U481 ( .A1(n87), .A2(n27), .Y(\ab[19][12] ) );
  AND2X1_RVT U482 ( .A1(n87), .A2(n25), .Y(\ab[19][11] ) );
  AND2X1_RVT U483 ( .A1(n87), .A2(n23), .Y(\ab[19][10] ) );
  AND2X1_RVT U484 ( .A1(n87), .A2(n3), .Y(\ab[19][0] ) );
  AND2X1_RVT U485 ( .A1(n85), .A2(n21), .Y(\ab[18][9] ) );
  AND2X1_RVT U486 ( .A1(n85), .A2(n19), .Y(\ab[18][8] ) );
  AND2X1_RVT U487 ( .A1(n85), .A2(n17), .Y(\ab[18][7] ) );
  AND2X1_RVT U488 ( .A1(n85), .A2(n15), .Y(\ab[18][6] ) );
  AND2X1_RVT U489 ( .A1(n85), .A2(n13), .Y(\ab[18][5] ) );
  AND2X1_RVT U490 ( .A1(n85), .A2(n11), .Y(\ab[18][4] ) );
  AND2X1_RVT U491 ( .A1(n85), .A2(n9), .Y(\ab[18][3] ) );
  AND2X1_RVT U492 ( .A1(n85), .A2(n7), .Y(\ab[18][2] ) );
  AND2X1_RVT U493 ( .A1(n85), .A2(n47), .Y(\ab[18][22] ) );
  AND2X1_RVT U494 ( .A1(n85), .A2(n45), .Y(\ab[18][21] ) );
  AND2X1_RVT U495 ( .A1(n85), .A2(n43), .Y(\ab[18][20] ) );
  AND2X1_RVT U496 ( .A1(n85), .A2(n5), .Y(\ab[18][1] ) );
  AND2X1_RVT U497 ( .A1(n85), .A2(n41), .Y(\ab[18][19] ) );
  AND2X1_RVT U498 ( .A1(n85), .A2(n39), .Y(\ab[18][18] ) );
  AND2X1_RVT U499 ( .A1(n85), .A2(n37), .Y(\ab[18][17] ) );
  AND2X1_RVT U500 ( .A1(n85), .A2(n35), .Y(\ab[18][16] ) );
  AND2X1_RVT U501 ( .A1(n85), .A2(n33), .Y(\ab[18][15] ) );
  AND2X1_RVT U502 ( .A1(n85), .A2(n31), .Y(\ab[18][14] ) );
  AND2X1_RVT U503 ( .A1(n85), .A2(n29), .Y(\ab[18][13] ) );
  AND2X1_RVT U504 ( .A1(n85), .A2(n27), .Y(\ab[18][12] ) );
  AND2X1_RVT U505 ( .A1(n85), .A2(n25), .Y(\ab[18][11] ) );
  AND2X1_RVT U506 ( .A1(n85), .A2(n23), .Y(\ab[18][10] ) );
  AND2X1_RVT U507 ( .A1(n85), .A2(n3), .Y(\ab[18][0] ) );
  AND2X1_RVT U508 ( .A1(n83), .A2(n21), .Y(\ab[17][9] ) );
  AND2X1_RVT U509 ( .A1(n83), .A2(n19), .Y(\ab[17][8] ) );
  AND2X1_RVT U510 ( .A1(n83), .A2(n17), .Y(\ab[17][7] ) );
  AND2X1_RVT U511 ( .A1(n83), .A2(n15), .Y(\ab[17][6] ) );
  AND2X1_RVT U512 ( .A1(n83), .A2(n13), .Y(\ab[17][5] ) );
  AND2X1_RVT U513 ( .A1(n83), .A2(n11), .Y(\ab[17][4] ) );
  AND2X1_RVT U514 ( .A1(n83), .A2(n9), .Y(\ab[17][3] ) );
  AND2X1_RVT U515 ( .A1(n83), .A2(n7), .Y(\ab[17][2] ) );
  AND2X1_RVT U516 ( .A1(n83), .A2(n47), .Y(\ab[17][22] ) );
  AND2X1_RVT U517 ( .A1(n83), .A2(n45), .Y(\ab[17][21] ) );
  AND2X1_RVT U518 ( .A1(n83), .A2(n43), .Y(\ab[17][20] ) );
  AND2X1_RVT U519 ( .A1(n83), .A2(n5), .Y(\ab[17][1] ) );
  AND2X1_RVT U520 ( .A1(n83), .A2(n41), .Y(\ab[17][19] ) );
  AND2X1_RVT U521 ( .A1(n83), .A2(n39), .Y(\ab[17][18] ) );
  AND2X1_RVT U522 ( .A1(n83), .A2(n37), .Y(\ab[17][17] ) );
  AND2X1_RVT U523 ( .A1(n83), .A2(n35), .Y(\ab[17][16] ) );
  AND2X1_RVT U524 ( .A1(n83), .A2(n33), .Y(\ab[17][15] ) );
  AND2X1_RVT U525 ( .A1(n83), .A2(n31), .Y(\ab[17][14] ) );
  AND2X1_RVT U526 ( .A1(n83), .A2(n29), .Y(\ab[17][13] ) );
  AND2X1_RVT U527 ( .A1(n83), .A2(n27), .Y(\ab[17][12] ) );
  AND2X1_RVT U528 ( .A1(n83), .A2(n25), .Y(\ab[17][11] ) );
  AND2X1_RVT U529 ( .A1(n83), .A2(n23), .Y(\ab[17][10] ) );
  AND2X1_RVT U530 ( .A1(n83), .A2(n3), .Y(\ab[17][0] ) );
  AND2X1_RVT U531 ( .A1(n81), .A2(n21), .Y(\ab[16][9] ) );
  AND2X1_RVT U532 ( .A1(n81), .A2(n19), .Y(\ab[16][8] ) );
  AND2X1_RVT U533 ( .A1(n81), .A2(n17), .Y(\ab[16][7] ) );
  AND2X1_RVT U534 ( .A1(n81), .A2(n15), .Y(\ab[16][6] ) );
  AND2X1_RVT U535 ( .A1(n81), .A2(n13), .Y(\ab[16][5] ) );
  AND2X1_RVT U536 ( .A1(n81), .A2(n11), .Y(\ab[16][4] ) );
  AND2X1_RVT U537 ( .A1(n81), .A2(n9), .Y(\ab[16][3] ) );
  AND2X1_RVT U538 ( .A1(n81), .A2(n7), .Y(\ab[16][2] ) );
  AND2X1_RVT U539 ( .A1(n81), .A2(n47), .Y(\ab[16][22] ) );
  AND2X1_RVT U540 ( .A1(n81), .A2(n45), .Y(\ab[16][21] ) );
  AND2X1_RVT U541 ( .A1(n81), .A2(n43), .Y(\ab[16][20] ) );
  AND2X1_RVT U542 ( .A1(n81), .A2(n5), .Y(\ab[16][1] ) );
  AND2X1_RVT U543 ( .A1(n81), .A2(n41), .Y(\ab[16][19] ) );
  AND2X1_RVT U544 ( .A1(n81), .A2(n39), .Y(\ab[16][18] ) );
  AND2X1_RVT U545 ( .A1(n81), .A2(n37), .Y(\ab[16][17] ) );
  AND2X1_RVT U546 ( .A1(n81), .A2(n35), .Y(\ab[16][16] ) );
  AND2X1_RVT U547 ( .A1(n81), .A2(n33), .Y(\ab[16][15] ) );
  AND2X1_RVT U548 ( .A1(n81), .A2(n31), .Y(\ab[16][14] ) );
  AND2X1_RVT U549 ( .A1(n81), .A2(n29), .Y(\ab[16][13] ) );
  AND2X1_RVT U550 ( .A1(n81), .A2(n27), .Y(\ab[16][12] ) );
  AND2X1_RVT U551 ( .A1(n81), .A2(n25), .Y(\ab[16][11] ) );
  AND2X1_RVT U552 ( .A1(n81), .A2(n23), .Y(\ab[16][10] ) );
  AND2X1_RVT U553 ( .A1(n81), .A2(n3), .Y(\ab[16][0] ) );
  AND2X1_RVT U554 ( .A1(n79), .A2(n21), .Y(\ab[15][9] ) );
  AND2X1_RVT U555 ( .A1(n79), .A2(n19), .Y(\ab[15][8] ) );
  AND2X1_RVT U556 ( .A1(n79), .A2(n17), .Y(\ab[15][7] ) );
  AND2X1_RVT U557 ( .A1(n79), .A2(n15), .Y(\ab[15][6] ) );
  AND2X1_RVT U558 ( .A1(n79), .A2(n13), .Y(\ab[15][5] ) );
  AND2X1_RVT U559 ( .A1(n79), .A2(n11), .Y(\ab[15][4] ) );
  AND2X1_RVT U560 ( .A1(n79), .A2(n9), .Y(\ab[15][3] ) );
  AND2X1_RVT U561 ( .A1(n79), .A2(n7), .Y(\ab[15][2] ) );
  AND2X1_RVT U562 ( .A1(n79), .A2(n47), .Y(\ab[15][22] ) );
  AND2X1_RVT U563 ( .A1(n79), .A2(n45), .Y(\ab[15][21] ) );
  AND2X1_RVT U564 ( .A1(n79), .A2(n43), .Y(\ab[15][20] ) );
  AND2X1_RVT U565 ( .A1(n79), .A2(n5), .Y(\ab[15][1] ) );
  AND2X1_RVT U566 ( .A1(n79), .A2(n41), .Y(\ab[15][19] ) );
  AND2X1_RVT U567 ( .A1(n79), .A2(n39), .Y(\ab[15][18] ) );
  AND2X1_RVT U568 ( .A1(n79), .A2(n37), .Y(\ab[15][17] ) );
  AND2X1_RVT U569 ( .A1(n79), .A2(n35), .Y(\ab[15][16] ) );
  AND2X1_RVT U570 ( .A1(n79), .A2(n33), .Y(\ab[15][15] ) );
  AND2X1_RVT U571 ( .A1(n79), .A2(n31), .Y(\ab[15][14] ) );
  AND2X1_RVT U572 ( .A1(n79), .A2(n29), .Y(\ab[15][13] ) );
  AND2X1_RVT U573 ( .A1(n79), .A2(n27), .Y(\ab[15][12] ) );
  AND2X1_RVT U574 ( .A1(n79), .A2(n25), .Y(\ab[15][11] ) );
  AND2X1_RVT U575 ( .A1(n79), .A2(n23), .Y(\ab[15][10] ) );
  AND2X1_RVT U576 ( .A1(n79), .A2(n3), .Y(\ab[15][0] ) );
  AND2X1_RVT U577 ( .A1(n77), .A2(n21), .Y(\ab[14][9] ) );
  AND2X1_RVT U578 ( .A1(n77), .A2(n19), .Y(\ab[14][8] ) );
  AND2X1_RVT U579 ( .A1(n77), .A2(n17), .Y(\ab[14][7] ) );
  AND2X1_RVT U580 ( .A1(n77), .A2(n15), .Y(\ab[14][6] ) );
  AND2X1_RVT U581 ( .A1(n77), .A2(n13), .Y(\ab[14][5] ) );
  AND2X1_RVT U582 ( .A1(n77), .A2(n11), .Y(\ab[14][4] ) );
  AND2X1_RVT U583 ( .A1(n77), .A2(n9), .Y(\ab[14][3] ) );
  AND2X1_RVT U584 ( .A1(n77), .A2(n7), .Y(\ab[14][2] ) );
  AND2X1_RVT U585 ( .A1(n77), .A2(n47), .Y(\ab[14][22] ) );
  AND2X1_RVT U586 ( .A1(n77), .A2(n45), .Y(\ab[14][21] ) );
  AND2X1_RVT U587 ( .A1(n77), .A2(n43), .Y(\ab[14][20] ) );
  AND2X1_RVT U588 ( .A1(n77), .A2(n5), .Y(\ab[14][1] ) );
  AND2X1_RVT U589 ( .A1(n77), .A2(n41), .Y(\ab[14][19] ) );
  AND2X1_RVT U590 ( .A1(n77), .A2(n39), .Y(\ab[14][18] ) );
  AND2X1_RVT U591 ( .A1(n77), .A2(n37), .Y(\ab[14][17] ) );
  AND2X1_RVT U592 ( .A1(n77), .A2(n35), .Y(\ab[14][16] ) );
  AND2X1_RVT U593 ( .A1(n77), .A2(n33), .Y(\ab[14][15] ) );
  AND2X1_RVT U594 ( .A1(n77), .A2(n31), .Y(\ab[14][14] ) );
  AND2X1_RVT U595 ( .A1(n77), .A2(n29), .Y(\ab[14][13] ) );
  AND2X1_RVT U596 ( .A1(n77), .A2(n27), .Y(\ab[14][12] ) );
  AND2X1_RVT U597 ( .A1(n77), .A2(n25), .Y(\ab[14][11] ) );
  AND2X1_RVT U598 ( .A1(n77), .A2(n23), .Y(\ab[14][10] ) );
  AND2X1_RVT U599 ( .A1(n77), .A2(n3), .Y(\ab[14][0] ) );
  AND2X1_RVT U600 ( .A1(n75), .A2(n21), .Y(\ab[13][9] ) );
  AND2X1_RVT U601 ( .A1(n75), .A2(n19), .Y(\ab[13][8] ) );
  AND2X1_RVT U602 ( .A1(n75), .A2(n17), .Y(\ab[13][7] ) );
  AND2X1_RVT U603 ( .A1(n75), .A2(n15), .Y(\ab[13][6] ) );
  AND2X1_RVT U604 ( .A1(n75), .A2(n13), .Y(\ab[13][5] ) );
  AND2X1_RVT U605 ( .A1(n75), .A2(n11), .Y(\ab[13][4] ) );
  AND2X1_RVT U606 ( .A1(n75), .A2(n9), .Y(\ab[13][3] ) );
  AND2X1_RVT U607 ( .A1(n75), .A2(n7), .Y(\ab[13][2] ) );
  AND2X1_RVT U608 ( .A1(n75), .A2(n47), .Y(\ab[13][22] ) );
  AND2X1_RVT U609 ( .A1(n75), .A2(n45), .Y(\ab[13][21] ) );
  AND2X1_RVT U610 ( .A1(n75), .A2(n43), .Y(\ab[13][20] ) );
  AND2X1_RVT U611 ( .A1(n75), .A2(n5), .Y(\ab[13][1] ) );
  AND2X1_RVT U612 ( .A1(n75), .A2(n41), .Y(\ab[13][19] ) );
  AND2X1_RVT U613 ( .A1(n75), .A2(n39), .Y(\ab[13][18] ) );
  AND2X1_RVT U614 ( .A1(n75), .A2(n37), .Y(\ab[13][17] ) );
  AND2X1_RVT U615 ( .A1(n75), .A2(n35), .Y(\ab[13][16] ) );
  AND2X1_RVT U616 ( .A1(n75), .A2(n33), .Y(\ab[13][15] ) );
  AND2X1_RVT U617 ( .A1(n75), .A2(n31), .Y(\ab[13][14] ) );
  AND2X1_RVT U618 ( .A1(n75), .A2(n29), .Y(\ab[13][13] ) );
  AND2X1_RVT U619 ( .A1(n75), .A2(n27), .Y(\ab[13][12] ) );
  AND2X1_RVT U620 ( .A1(n75), .A2(n25), .Y(\ab[13][11] ) );
  AND2X1_RVT U621 ( .A1(n75), .A2(n23), .Y(\ab[13][10] ) );
  AND2X1_RVT U622 ( .A1(n75), .A2(n3), .Y(\ab[13][0] ) );
  AND2X1_RVT U623 ( .A1(n73), .A2(n21), .Y(\ab[12][9] ) );
  AND2X1_RVT U624 ( .A1(n73), .A2(n19), .Y(\ab[12][8] ) );
  AND2X1_RVT U625 ( .A1(n73), .A2(n17), .Y(\ab[12][7] ) );
  AND2X1_RVT U626 ( .A1(n73), .A2(n15), .Y(\ab[12][6] ) );
  AND2X1_RVT U627 ( .A1(n73), .A2(n13), .Y(\ab[12][5] ) );
  AND2X1_RVT U628 ( .A1(n73), .A2(n11), .Y(\ab[12][4] ) );
  AND2X1_RVT U629 ( .A1(n73), .A2(n9), .Y(\ab[12][3] ) );
  AND2X1_RVT U630 ( .A1(n73), .A2(n7), .Y(\ab[12][2] ) );
  AND2X1_RVT U631 ( .A1(n73), .A2(n47), .Y(\ab[12][22] ) );
  AND2X1_RVT U632 ( .A1(n73), .A2(n45), .Y(\ab[12][21] ) );
  AND2X1_RVT U633 ( .A1(n73), .A2(n43), .Y(\ab[12][20] ) );
  AND2X1_RVT U634 ( .A1(n73), .A2(n5), .Y(\ab[12][1] ) );
  AND2X1_RVT U635 ( .A1(n73), .A2(n41), .Y(\ab[12][19] ) );
  AND2X1_RVT U636 ( .A1(n73), .A2(n39), .Y(\ab[12][18] ) );
  AND2X1_RVT U637 ( .A1(n73), .A2(n37), .Y(\ab[12][17] ) );
  AND2X1_RVT U638 ( .A1(n73), .A2(n35), .Y(\ab[12][16] ) );
  AND2X1_RVT U639 ( .A1(n73), .A2(n33), .Y(\ab[12][15] ) );
  AND2X1_RVT U640 ( .A1(n73), .A2(n31), .Y(\ab[12][14] ) );
  AND2X1_RVT U641 ( .A1(n73), .A2(n29), .Y(\ab[12][13] ) );
  AND2X1_RVT U642 ( .A1(n73), .A2(n27), .Y(\ab[12][12] ) );
  AND2X1_RVT U643 ( .A1(n73), .A2(n25), .Y(\ab[12][11] ) );
  AND2X1_RVT U644 ( .A1(n73), .A2(n23), .Y(\ab[12][10] ) );
  AND2X1_RVT U645 ( .A1(n73), .A2(n3), .Y(\ab[12][0] ) );
  AND2X1_RVT U646 ( .A1(n71), .A2(n21), .Y(\ab[11][9] ) );
  AND2X1_RVT U647 ( .A1(n71), .A2(n19), .Y(\ab[11][8] ) );
  AND2X1_RVT U648 ( .A1(n71), .A2(n17), .Y(\ab[11][7] ) );
  AND2X1_RVT U649 ( .A1(n71), .A2(n15), .Y(\ab[11][6] ) );
  AND2X1_RVT U650 ( .A1(n71), .A2(n13), .Y(\ab[11][5] ) );
  AND2X1_RVT U651 ( .A1(n71), .A2(n11), .Y(\ab[11][4] ) );
  AND2X1_RVT U652 ( .A1(n71), .A2(n9), .Y(\ab[11][3] ) );
  AND2X1_RVT U653 ( .A1(n71), .A2(n7), .Y(\ab[11][2] ) );
  AND2X1_RVT U654 ( .A1(n71), .A2(n47), .Y(\ab[11][22] ) );
  AND2X1_RVT U655 ( .A1(n71), .A2(n45), .Y(\ab[11][21] ) );
  AND2X1_RVT U656 ( .A1(n71), .A2(n43), .Y(\ab[11][20] ) );
  AND2X1_RVT U657 ( .A1(n71), .A2(n5), .Y(\ab[11][1] ) );
  AND2X1_RVT U658 ( .A1(n71), .A2(n41), .Y(\ab[11][19] ) );
  AND2X1_RVT U659 ( .A1(n71), .A2(n39), .Y(\ab[11][18] ) );
  AND2X1_RVT U660 ( .A1(n71), .A2(n37), .Y(\ab[11][17] ) );
  AND2X1_RVT U661 ( .A1(n71), .A2(n35), .Y(\ab[11][16] ) );
  AND2X1_RVT U662 ( .A1(n71), .A2(n33), .Y(\ab[11][15] ) );
  AND2X1_RVT U663 ( .A1(n71), .A2(n31), .Y(\ab[11][14] ) );
  AND2X1_RVT U664 ( .A1(n71), .A2(n29), .Y(\ab[11][13] ) );
  AND2X1_RVT U665 ( .A1(n71), .A2(n27), .Y(\ab[11][12] ) );
  AND2X1_RVT U666 ( .A1(n71), .A2(n25), .Y(\ab[11][11] ) );
  AND2X1_RVT U667 ( .A1(n71), .A2(n23), .Y(\ab[11][10] ) );
  AND2X1_RVT U668 ( .A1(n71), .A2(n3), .Y(\ab[11][0] ) );
  AND2X1_RVT U669 ( .A1(n69), .A2(n21), .Y(\ab[10][9] ) );
  AND2X1_RVT U670 ( .A1(n69), .A2(n19), .Y(\ab[10][8] ) );
  AND2X1_RVT U671 ( .A1(n69), .A2(n17), .Y(\ab[10][7] ) );
  AND2X1_RVT U672 ( .A1(n69), .A2(n15), .Y(\ab[10][6] ) );
  AND2X1_RVT U673 ( .A1(n69), .A2(n13), .Y(\ab[10][5] ) );
  AND2X1_RVT U674 ( .A1(n69), .A2(n11), .Y(\ab[10][4] ) );
  AND2X1_RVT U675 ( .A1(n69), .A2(n9), .Y(\ab[10][3] ) );
  AND2X1_RVT U676 ( .A1(n69), .A2(n7), .Y(\ab[10][2] ) );
  AND2X1_RVT U677 ( .A1(n69), .A2(n47), .Y(\ab[10][22] ) );
  AND2X1_RVT U678 ( .A1(n69), .A2(n45), .Y(\ab[10][21] ) );
  AND2X1_RVT U679 ( .A1(n69), .A2(n43), .Y(\ab[10][20] ) );
  AND2X1_RVT U680 ( .A1(n69), .A2(n5), .Y(\ab[10][1] ) );
  AND2X1_RVT U681 ( .A1(n69), .A2(n41), .Y(\ab[10][19] ) );
  AND2X1_RVT U682 ( .A1(n69), .A2(n39), .Y(\ab[10][18] ) );
  AND2X1_RVT U683 ( .A1(n69), .A2(n37), .Y(\ab[10][17] ) );
  AND2X1_RVT U684 ( .A1(n69), .A2(n35), .Y(\ab[10][16] ) );
  AND2X1_RVT U685 ( .A1(n69), .A2(n33), .Y(\ab[10][15] ) );
  AND2X1_RVT U686 ( .A1(n69), .A2(n31), .Y(\ab[10][14] ) );
  AND2X1_RVT U687 ( .A1(n69), .A2(n29), .Y(\ab[10][13] ) );
  AND2X1_RVT U688 ( .A1(n69), .A2(n27), .Y(\ab[10][12] ) );
  AND2X1_RVT U689 ( .A1(n69), .A2(n25), .Y(\ab[10][11] ) );
  AND2X1_RVT U690 ( .A1(n69), .A2(n23), .Y(\ab[10][10] ) );
  AND2X1_RVT U691 ( .A1(n69), .A2(n3), .Y(\ab[10][0] ) );
  AND2X1_RVT U692 ( .A1(n49), .A2(n21), .Y(\ab[0][9] ) );
  AND2X1_RVT U693 ( .A1(n49), .A2(n19), .Y(\ab[0][8] ) );
  AND2X1_RVT U694 ( .A1(n49), .A2(n17), .Y(\ab[0][7] ) );
  AND2X1_RVT U695 ( .A1(n49), .A2(n15), .Y(\ab[0][6] ) );
  AND2X1_RVT U696 ( .A1(n49), .A2(n13), .Y(\ab[0][5] ) );
  AND2X1_RVT U697 ( .A1(n49), .A2(n11), .Y(\ab[0][4] ) );
  AND2X1_RVT U698 ( .A1(n49), .A2(n9), .Y(\ab[0][3] ) );
  AND2X1_RVT U699 ( .A1(n49), .A2(n7), .Y(\ab[0][2] ) );
  AND2X1_RVT U700 ( .A1(n49), .A2(n47), .Y(\ab[0][22] ) );
  AND2X1_RVT U701 ( .A1(n49), .A2(n45), .Y(\ab[0][21] ) );
  AND2X1_RVT U702 ( .A1(n49), .A2(n43), .Y(\ab[0][20] ) );
  AND2X1_RVT U703 ( .A1(n49), .A2(n5), .Y(\ab[0][1] ) );
  AND2X1_RVT U704 ( .A1(n49), .A2(n41), .Y(\ab[0][19] ) );
  AND2X1_RVT U705 ( .A1(n49), .A2(n39), .Y(\ab[0][18] ) );
  AND2X1_RVT U706 ( .A1(n49), .A2(n37), .Y(\ab[0][17] ) );
  AND2X1_RVT U707 ( .A1(n49), .A2(n35), .Y(\ab[0][16] ) );
  AND2X1_RVT U708 ( .A1(n49), .A2(n33), .Y(\ab[0][15] ) );
  AND2X1_RVT U709 ( .A1(n49), .A2(n31), .Y(\ab[0][14] ) );
  AND2X1_RVT U710 ( .A1(n49), .A2(n29), .Y(\ab[0][13] ) );
  AND2X1_RVT U711 ( .A1(n49), .A2(n27), .Y(\ab[0][12] ) );
  AND2X1_RVT U712 ( .A1(n49), .A2(n25), .Y(\ab[0][11] ) );
  AND2X1_RVT U713 ( .A1(n49), .A2(n23), .Y(\ab[0][10] ) );
  AND2X1_RVT U714 ( .A1(n49), .A2(n3), .Y(PRODUCT[0]) );
endmodule


module FPU_CAL_DW01_add_3 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  XOR2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
  XOR2X1_RVT U2 ( .A1(B[8]), .A2(carry[8]), .Y(SUM[8]) );
  AND2X1_RVT U3 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
endmodule


module FPU_CAL_DW01_inc_4 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1_RVT U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1_RVT U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1_RVT U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1_RVT U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1_RVT U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1_RVT U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1_RVT U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0_RVT U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1_RVT U2 ( .A1(carry[8]), .A2(A[8]), .Y(SUM[8]) );
endmodule


module FPU_CAL_DW_div_uns_2 ( a, b, quotient, remainder, divide_by_0 );
  input [47:0] a;
  input [23:0] b;
  output [47:0] quotient;
  output [23:0] remainder;
  output divide_by_0;
  wire   n629, \u_div/SumTmp[15][1] , \u_div/SumTmp[15][2] ,
         \u_div/SumTmp[15][3] , \u_div/SumTmp[15][4] , \u_div/SumTmp[15][5] ,
         \u_div/SumTmp[15][6] , \u_div/SumTmp[15][7] , \u_div/SumTmp[15][8] ,
         \u_div/SumTmp[15][9] , \u_div/SumTmp[15][10] , \u_div/SumTmp[15][11] ,
         \u_div/SumTmp[15][12] , \u_div/SumTmp[15][13] ,
         \u_div/SumTmp[15][14] , \u_div/SumTmp[15][15] ,
         \u_div/SumTmp[15][16] , \u_div/SumTmp[15][17] ,
         \u_div/SumTmp[15][18] , \u_div/SumTmp[15][19] ,
         \u_div/SumTmp[15][20] , \u_div/SumTmp[15][21] ,
         \u_div/SumTmp[15][22] , \u_div/SumTmp[15][23] , \u_div/SumTmp[16][1] ,
         \u_div/SumTmp[16][2] , \u_div/SumTmp[16][3] , \u_div/SumTmp[16][4] ,
         \u_div/SumTmp[16][5] , \u_div/SumTmp[16][6] , \u_div/SumTmp[16][7] ,
         \u_div/SumTmp[16][8] , \u_div/SumTmp[16][9] , \u_div/SumTmp[16][10] ,
         \u_div/SumTmp[16][11] , \u_div/SumTmp[16][12] ,
         \u_div/SumTmp[16][13] , \u_div/SumTmp[16][14] ,
         \u_div/SumTmp[16][15] , \u_div/SumTmp[16][16] ,
         \u_div/SumTmp[16][17] , \u_div/SumTmp[16][18] ,
         \u_div/SumTmp[16][19] , \u_div/SumTmp[16][20] ,
         \u_div/SumTmp[16][21] , \u_div/SumTmp[16][22] ,
         \u_div/SumTmp[16][23] , \u_div/SumTmp[17][1] , \u_div/SumTmp[17][2] ,
         \u_div/SumTmp[17][3] , \u_div/SumTmp[17][4] , \u_div/SumTmp[17][5] ,
         \u_div/SumTmp[17][6] , \u_div/SumTmp[17][7] , \u_div/SumTmp[17][8] ,
         \u_div/SumTmp[17][9] , \u_div/SumTmp[17][10] , \u_div/SumTmp[17][11] ,
         \u_div/SumTmp[17][12] , \u_div/SumTmp[17][13] ,
         \u_div/SumTmp[17][14] , \u_div/SumTmp[17][15] ,
         \u_div/SumTmp[17][16] , \u_div/SumTmp[17][17] ,
         \u_div/SumTmp[17][18] , \u_div/SumTmp[17][19] ,
         \u_div/SumTmp[17][20] , \u_div/SumTmp[17][21] ,
         \u_div/SumTmp[17][22] , \u_div/SumTmp[17][23] , \u_div/SumTmp[18][0] ,
         \u_div/SumTmp[18][1] , \u_div/SumTmp[18][2] , \u_div/SumTmp[18][3] ,
         \u_div/SumTmp[18][4] , \u_div/SumTmp[18][5] , \u_div/SumTmp[18][6] ,
         \u_div/SumTmp[18][7] , \u_div/SumTmp[18][8] , \u_div/SumTmp[18][9] ,
         \u_div/SumTmp[18][10] , \u_div/SumTmp[18][11] ,
         \u_div/SumTmp[18][12] , \u_div/SumTmp[18][13] ,
         \u_div/SumTmp[18][14] , \u_div/SumTmp[18][15] ,
         \u_div/SumTmp[18][16] , \u_div/SumTmp[18][17] ,
         \u_div/SumTmp[18][18] , \u_div/SumTmp[18][19] ,
         \u_div/SumTmp[18][20] , \u_div/SumTmp[18][21] ,
         \u_div/SumTmp[18][22] , \u_div/SumTmp[18][23] , \u_div/SumTmp[19][0] ,
         \u_div/SumTmp[19][1] , \u_div/SumTmp[19][2] , \u_div/SumTmp[19][3] ,
         \u_div/SumTmp[19][4] , \u_div/SumTmp[19][5] , \u_div/SumTmp[19][6] ,
         \u_div/SumTmp[19][7] , \u_div/SumTmp[19][8] , \u_div/SumTmp[19][9] ,
         \u_div/SumTmp[19][11] , \u_div/SumTmp[19][12] ,
         \u_div/SumTmp[19][13] , \u_div/SumTmp[19][14] ,
         \u_div/SumTmp[19][15] , \u_div/SumTmp[19][16] ,
         \u_div/SumTmp[19][17] , \u_div/SumTmp[19][18] ,
         \u_div/SumTmp[19][19] , \u_div/SumTmp[19][20] ,
         \u_div/SumTmp[19][21] , \u_div/SumTmp[19][22] ,
         \u_div/SumTmp[19][23] , \u_div/SumTmp[20][0] , \u_div/SumTmp[20][1] ,
         \u_div/SumTmp[20][2] , \u_div/SumTmp[20][3] , \u_div/SumTmp[20][4] ,
         \u_div/SumTmp[20][5] , \u_div/SumTmp[20][6] , \u_div/SumTmp[20][7] ,
         \u_div/SumTmp[20][8] , \u_div/SumTmp[20][9] , \u_div/SumTmp[20][10] ,
         \u_div/SumTmp[20][11] , \u_div/SumTmp[20][12] ,
         \u_div/SumTmp[20][13] , \u_div/SumTmp[20][14] ,
         \u_div/SumTmp[20][15] , \u_div/SumTmp[20][16] ,
         \u_div/SumTmp[20][17] , \u_div/SumTmp[20][18] ,
         \u_div/SumTmp[20][19] , \u_div/SumTmp[20][20] ,
         \u_div/SumTmp[20][21] , \u_div/SumTmp[20][22] ,
         \u_div/SumTmp[20][23] , \u_div/SumTmp[21][0] , \u_div/SumTmp[21][1] ,
         \u_div/SumTmp[21][2] , \u_div/SumTmp[21][3] , \u_div/SumTmp[21][4] ,
         \u_div/SumTmp[21][5] , \u_div/SumTmp[21][6] , \u_div/SumTmp[21][7] ,
         \u_div/SumTmp[21][8] , \u_div/SumTmp[21][9] , \u_div/SumTmp[21][10] ,
         \u_div/SumTmp[21][11] , \u_div/SumTmp[21][12] ,
         \u_div/SumTmp[21][13] , \u_div/SumTmp[21][14] ,
         \u_div/SumTmp[21][15] , \u_div/SumTmp[21][16] ,
         \u_div/SumTmp[21][17] , \u_div/SumTmp[21][18] ,
         \u_div/SumTmp[21][19] , \u_div/SumTmp[21][20] ,
         \u_div/SumTmp[21][21] , \u_div/SumTmp[21][22] ,
         \u_div/SumTmp[21][23] , \u_div/SumTmp[22][0] , \u_div/SumTmp[22][1] ,
         \u_div/SumTmp[22][2] , \u_div/SumTmp[22][3] , \u_div/SumTmp[22][4] ,
         \u_div/SumTmp[22][5] , \u_div/SumTmp[22][6] , \u_div/SumTmp[22][7] ,
         \u_div/SumTmp[22][8] , \u_div/SumTmp[22][9] , \u_div/SumTmp[22][10] ,
         \u_div/SumTmp[22][11] , \u_div/SumTmp[22][12] ,
         \u_div/SumTmp[22][13] , \u_div/SumTmp[22][14] ,
         \u_div/SumTmp[22][15] , \u_div/SumTmp[22][16] ,
         \u_div/SumTmp[22][17] , \u_div/SumTmp[22][18] ,
         \u_div/SumTmp[22][19] , \u_div/SumTmp[22][20] ,
         \u_div/SumTmp[22][21] , \u_div/SumTmp[22][22] ,
         \u_div/SumTmp[22][23] , \u_div/SumTmp[23][0] , \u_div/SumTmp[23][1] ,
         \u_div/SumTmp[23][2] , \u_div/SumTmp[23][3] , \u_div/SumTmp[23][4] ,
         \u_div/SumTmp[23][5] , \u_div/SumTmp[23][6] , \u_div/SumTmp[23][7] ,
         \u_div/SumTmp[23][8] , \u_div/SumTmp[23][9] , \u_div/SumTmp[23][10] ,
         \u_div/SumTmp[23][11] , \u_div/SumTmp[23][12] ,
         \u_div/SumTmp[23][13] , \u_div/SumTmp[23][14] ,
         \u_div/SumTmp[23][15] , \u_div/SumTmp[23][16] ,
         \u_div/SumTmp[23][17] , \u_div/SumTmp[23][18] ,
         \u_div/SumTmp[23][19] , \u_div/SumTmp[23][20] ,
         \u_div/SumTmp[23][21] , \u_div/SumTmp[23][22] ,
         \u_div/SumTmp[23][23] , \u_div/SumTmp[24][1] , \u_div/SumTmp[24][2] ,
         \u_div/SumTmp[24][3] , \u_div/SumTmp[24][4] , \u_div/SumTmp[24][5] ,
         \u_div/SumTmp[24][6] , \u_div/SumTmp[24][7] , \u_div/SumTmp[24][8] ,
         \u_div/SumTmp[24][9] , \u_div/SumTmp[24][10] , \u_div/SumTmp[24][11] ,
         \u_div/SumTmp[24][12] , \u_div/SumTmp[24][13] ,
         \u_div/SumTmp[24][14] , \u_div/SumTmp[24][15] ,
         \u_div/SumTmp[24][16] , \u_div/SumTmp[24][17] ,
         \u_div/SumTmp[24][18] , \u_div/SumTmp[24][19] ,
         \u_div/SumTmp[24][20] , \u_div/SumTmp[24][21] ,
         \u_div/SumTmp[24][22] , \u_div/SumTmp[24][23] , \u_div/CryTmp[14][2] ,
         \u_div/CryTmp[14][3] , \u_div/CryTmp[14][4] , \u_div/CryTmp[14][5] ,
         \u_div/CryTmp[14][6] , \u_div/CryTmp[14][7] , \u_div/CryTmp[14][8] ,
         \u_div/CryTmp[14][9] , \u_div/CryTmp[14][10] , \u_div/CryTmp[14][11] ,
         \u_div/CryTmp[14][12] , \u_div/CryTmp[14][13] ,
         \u_div/CryTmp[14][14] , \u_div/CryTmp[14][15] ,
         \u_div/CryTmp[14][16] , \u_div/CryTmp[14][17] ,
         \u_div/CryTmp[14][18] , \u_div/CryTmp[14][19] ,
         \u_div/CryTmp[14][20] , \u_div/CryTmp[14][21] ,
         \u_div/CryTmp[14][22] , \u_div/CryTmp[14][23] ,
         \u_div/CryTmp[14][24] , \u_div/CryTmp[15][2] , \u_div/CryTmp[15][3] ,
         \u_div/CryTmp[15][4] , \u_div/CryTmp[15][5] , \u_div/CryTmp[15][6] ,
         \u_div/CryTmp[15][7] , \u_div/CryTmp[15][8] , \u_div/CryTmp[15][9] ,
         \u_div/CryTmp[15][10] , \u_div/CryTmp[15][11] ,
         \u_div/CryTmp[15][12] , \u_div/CryTmp[15][13] ,
         \u_div/CryTmp[15][14] , \u_div/CryTmp[15][15] ,
         \u_div/CryTmp[15][16] , \u_div/CryTmp[15][17] ,
         \u_div/CryTmp[15][18] , \u_div/CryTmp[15][19] ,
         \u_div/CryTmp[15][20] , \u_div/CryTmp[15][21] ,
         \u_div/CryTmp[15][22] , \u_div/CryTmp[15][23] ,
         \u_div/CryTmp[15][24] , \u_div/CryTmp[16][2] , \u_div/CryTmp[16][3] ,
         \u_div/CryTmp[16][4] , \u_div/CryTmp[16][5] , \u_div/CryTmp[16][6] ,
         \u_div/CryTmp[16][7] , \u_div/CryTmp[16][8] , \u_div/CryTmp[16][9] ,
         \u_div/CryTmp[16][10] , \u_div/CryTmp[16][11] ,
         \u_div/CryTmp[16][12] , \u_div/CryTmp[16][13] ,
         \u_div/CryTmp[16][14] , \u_div/CryTmp[16][15] ,
         \u_div/CryTmp[16][16] , \u_div/CryTmp[16][17] ,
         \u_div/CryTmp[16][18] , \u_div/CryTmp[16][19] ,
         \u_div/CryTmp[16][20] , \u_div/CryTmp[16][21] ,
         \u_div/CryTmp[16][22] , \u_div/CryTmp[16][23] ,
         \u_div/CryTmp[16][24] , \u_div/CryTmp[17][2] , \u_div/CryTmp[17][3] ,
         \u_div/CryTmp[17][4] , \u_div/CryTmp[17][5] , \u_div/CryTmp[17][6] ,
         \u_div/CryTmp[17][7] , \u_div/CryTmp[17][8] , \u_div/CryTmp[17][9] ,
         \u_div/CryTmp[17][10] , \u_div/CryTmp[17][11] ,
         \u_div/CryTmp[17][12] , \u_div/CryTmp[17][13] ,
         \u_div/CryTmp[17][14] , \u_div/CryTmp[17][15] ,
         \u_div/CryTmp[17][16] , \u_div/CryTmp[17][17] ,
         \u_div/CryTmp[17][18] , \u_div/CryTmp[17][19] ,
         \u_div/CryTmp[17][20] , \u_div/CryTmp[17][21] ,
         \u_div/CryTmp[17][22] , \u_div/CryTmp[17][23] ,
         \u_div/CryTmp[17][24] , \u_div/CryTmp[18][2] , \u_div/CryTmp[18][3] ,
         \u_div/CryTmp[18][4] , \u_div/CryTmp[18][5] , \u_div/CryTmp[18][6] ,
         \u_div/CryTmp[18][7] , \u_div/CryTmp[18][8] , \u_div/CryTmp[18][9] ,
         \u_div/CryTmp[18][10] , \u_div/CryTmp[18][11] ,
         \u_div/CryTmp[18][12] , \u_div/CryTmp[18][13] ,
         \u_div/CryTmp[18][14] , \u_div/CryTmp[18][15] ,
         \u_div/CryTmp[18][16] , \u_div/CryTmp[18][17] ,
         \u_div/CryTmp[18][18] , \u_div/CryTmp[18][19] ,
         \u_div/CryTmp[18][20] , \u_div/CryTmp[18][21] ,
         \u_div/CryTmp[18][22] , \u_div/CryTmp[18][23] ,
         \u_div/CryTmp[18][24] , \u_div/CryTmp[19][2] , \u_div/CryTmp[19][3] ,
         \u_div/CryTmp[19][4] , \u_div/CryTmp[19][5] , \u_div/CryTmp[19][6] ,
         \u_div/CryTmp[19][7] , \u_div/CryTmp[19][8] , \u_div/CryTmp[19][9] ,
         \u_div/CryTmp[19][10] , \u_div/CryTmp[19][11] ,
         \u_div/CryTmp[19][12] , \u_div/CryTmp[19][13] ,
         \u_div/CryTmp[19][14] , \u_div/CryTmp[19][15] ,
         \u_div/CryTmp[19][16] , \u_div/CryTmp[19][17] ,
         \u_div/CryTmp[19][18] , \u_div/CryTmp[19][19] ,
         \u_div/CryTmp[19][20] , \u_div/CryTmp[19][21] ,
         \u_div/CryTmp[19][22] , \u_div/CryTmp[19][23] ,
         \u_div/CryTmp[19][24] , \u_div/CryTmp[20][2] , \u_div/CryTmp[20][3] ,
         \u_div/CryTmp[20][4] , \u_div/CryTmp[20][5] , \u_div/CryTmp[20][6] ,
         \u_div/CryTmp[20][7] , \u_div/CryTmp[20][8] , \u_div/CryTmp[20][9] ,
         \u_div/CryTmp[20][10] , \u_div/CryTmp[20][11] ,
         \u_div/CryTmp[20][12] , \u_div/CryTmp[20][13] ,
         \u_div/CryTmp[20][14] , \u_div/CryTmp[20][15] ,
         \u_div/CryTmp[20][16] , \u_div/CryTmp[20][17] ,
         \u_div/CryTmp[20][18] , \u_div/CryTmp[20][19] ,
         \u_div/CryTmp[20][20] , \u_div/CryTmp[20][21] ,
         \u_div/CryTmp[20][22] , \u_div/CryTmp[20][23] , \u_div/CryTmp[21][2] ,
         \u_div/CryTmp[21][3] , \u_div/CryTmp[21][4] , \u_div/CryTmp[21][5] ,
         \u_div/CryTmp[21][6] , \u_div/CryTmp[21][7] , \u_div/CryTmp[21][8] ,
         \u_div/CryTmp[21][9] , \u_div/CryTmp[21][10] , \u_div/CryTmp[21][11] ,
         \u_div/CryTmp[21][12] , \u_div/CryTmp[21][13] ,
         \u_div/CryTmp[21][14] , \u_div/CryTmp[21][15] ,
         \u_div/CryTmp[21][16] , \u_div/CryTmp[21][17] ,
         \u_div/CryTmp[21][18] , \u_div/CryTmp[21][19] ,
         \u_div/CryTmp[21][20] , \u_div/CryTmp[21][21] ,
         \u_div/CryTmp[21][22] , \u_div/CryTmp[21][23] ,
         \u_div/CryTmp[21][24] , \u_div/CryTmp[22][2] , \u_div/CryTmp[22][3] ,
         \u_div/CryTmp[22][4] , \u_div/CryTmp[22][5] , \u_div/CryTmp[22][6] ,
         \u_div/CryTmp[22][7] , \u_div/CryTmp[22][8] , \u_div/CryTmp[22][9] ,
         \u_div/CryTmp[22][10] , \u_div/CryTmp[22][11] ,
         \u_div/CryTmp[22][12] , \u_div/CryTmp[22][13] ,
         \u_div/CryTmp[22][14] , \u_div/CryTmp[22][15] ,
         \u_div/CryTmp[22][16] , \u_div/CryTmp[22][17] ,
         \u_div/CryTmp[22][18] , \u_div/CryTmp[22][19] ,
         \u_div/CryTmp[22][20] , \u_div/CryTmp[22][21] ,
         \u_div/CryTmp[22][22] , \u_div/CryTmp[22][23] ,
         \u_div/CryTmp[22][24] , \u_div/CryTmp[23][1] , \u_div/CryTmp[23][2] ,
         \u_div/CryTmp[23][3] , \u_div/CryTmp[23][4] , \u_div/CryTmp[23][5] ,
         \u_div/CryTmp[23][6] , \u_div/CryTmp[23][7] , \u_div/CryTmp[23][8] ,
         \u_div/CryTmp[23][9] , \u_div/CryTmp[23][10] , \u_div/CryTmp[23][11] ,
         \u_div/CryTmp[23][12] , \u_div/CryTmp[23][13] ,
         \u_div/CryTmp[23][14] , \u_div/CryTmp[23][15] ,
         \u_div/CryTmp[23][16] , \u_div/CryTmp[23][17] ,
         \u_div/CryTmp[23][18] , \u_div/CryTmp[23][19] ,
         \u_div/CryTmp[23][20] , \u_div/CryTmp[23][21] ,
         \u_div/CryTmp[23][22] , \u_div/CryTmp[23][23] ,
         \u_div/CryTmp[23][24] , \u_div/CryTmp[24][1] , \u_div/CryTmp[24][2] ,
         \u_div/CryTmp[24][3] , \u_div/CryTmp[24][4] , \u_div/CryTmp[24][5] ,
         \u_div/CryTmp[24][6] , \u_div/CryTmp[24][7] , \u_div/CryTmp[24][8] ,
         \u_div/CryTmp[24][9] , \u_div/CryTmp[24][10] , \u_div/CryTmp[24][11] ,
         \u_div/CryTmp[24][12] , \u_div/CryTmp[24][13] ,
         \u_div/CryTmp[24][14] , \u_div/CryTmp[24][15] ,
         \u_div/CryTmp[24][16] , \u_div/CryTmp[24][17] ,
         \u_div/CryTmp[24][18] , \u_div/CryTmp[24][19] ,
         \u_div/CryTmp[24][20] , \u_div/CryTmp[24][21] ,
         \u_div/CryTmp[24][22] , \u_div/CryTmp[24][24] ,
         \u_div/PartRem[15][2] , \u_div/PartRem[15][3] ,
         \u_div/PartRem[15][4] , \u_div/PartRem[15][5] ,
         \u_div/PartRem[15][6] , \u_div/PartRem[15][7] ,
         \u_div/PartRem[15][8] , \u_div/PartRem[15][9] ,
         \u_div/PartRem[15][10] , \u_div/PartRem[15][11] ,
         \u_div/PartRem[15][12] , \u_div/PartRem[15][13] ,
         \u_div/PartRem[15][14] , \u_div/PartRem[15][15] ,
         \u_div/PartRem[15][16] , \u_div/PartRem[15][17] ,
         \u_div/PartRem[15][18] , \u_div/PartRem[15][19] ,
         \u_div/PartRem[15][20] , \u_div/PartRem[15][21] ,
         \u_div/PartRem[15][22] , \u_div/PartRem[15][23] ,
         \u_div/PartRem[15][24] , \u_div/PartRem[16][1] ,
         \u_div/PartRem[16][2] , \u_div/PartRem[16][3] ,
         \u_div/PartRem[16][4] , \u_div/PartRem[16][5] ,
         \u_div/PartRem[16][6] , \u_div/PartRem[16][7] ,
         \u_div/PartRem[16][8] , \u_div/PartRem[16][9] ,
         \u_div/PartRem[16][10] , \u_div/PartRem[16][11] ,
         \u_div/PartRem[16][12] , \u_div/PartRem[16][13] ,
         \u_div/PartRem[16][14] , \u_div/PartRem[16][15] ,
         \u_div/PartRem[16][16] , \u_div/PartRem[16][17] ,
         \u_div/PartRem[16][18] , \u_div/PartRem[16][19] ,
         \u_div/PartRem[16][20] , \u_div/PartRem[16][21] ,
         \u_div/PartRem[16][22] , \u_div/PartRem[16][23] ,
         \u_div/PartRem[16][24] , \u_div/PartRem[17][1] ,
         \u_div/PartRem[17][2] , \u_div/PartRem[17][3] ,
         \u_div/PartRem[17][4] , \u_div/PartRem[17][5] ,
         \u_div/PartRem[17][6] , \u_div/PartRem[17][7] ,
         \u_div/PartRem[17][8] , \u_div/PartRem[17][9] ,
         \u_div/PartRem[17][10] , \u_div/PartRem[17][11] ,
         \u_div/PartRem[17][12] , \u_div/PartRem[17][13] ,
         \u_div/PartRem[17][14] , \u_div/PartRem[17][15] ,
         \u_div/PartRem[17][16] , \u_div/PartRem[17][17] ,
         \u_div/PartRem[17][18] , \u_div/PartRem[17][19] ,
         \u_div/PartRem[17][20] , \u_div/PartRem[17][21] ,
         \u_div/PartRem[17][22] , \u_div/PartRem[17][23] ,
         \u_div/PartRem[17][24] , \u_div/PartRem[18][1] ,
         \u_div/PartRem[18][2] , \u_div/PartRem[18][3] ,
         \u_div/PartRem[18][4] , \u_div/PartRem[18][5] ,
         \u_div/PartRem[18][6] , \u_div/PartRem[18][7] ,
         \u_div/PartRem[18][8] , \u_div/PartRem[18][9] ,
         \u_div/PartRem[18][10] , \u_div/PartRem[18][11] ,
         \u_div/PartRem[18][12] , \u_div/PartRem[18][13] ,
         \u_div/PartRem[18][14] , \u_div/PartRem[18][15] ,
         \u_div/PartRem[18][16] , \u_div/PartRem[18][17] ,
         \u_div/PartRem[18][18] , \u_div/PartRem[18][19] ,
         \u_div/PartRem[18][20] , \u_div/PartRem[18][21] ,
         \u_div/PartRem[18][22] , \u_div/PartRem[18][23] ,
         \u_div/PartRem[18][24] , \u_div/PartRem[19][1] ,
         \u_div/PartRem[19][2] , \u_div/PartRem[19][3] ,
         \u_div/PartRem[19][4] , \u_div/PartRem[19][5] ,
         \u_div/PartRem[19][6] , \u_div/PartRem[19][7] ,
         \u_div/PartRem[19][8] , \u_div/PartRem[19][9] ,
         \u_div/PartRem[19][10] , \u_div/PartRem[19][11] ,
         \u_div/PartRem[19][12] , \u_div/PartRem[19][13] ,
         \u_div/PartRem[19][14] , \u_div/PartRem[19][15] ,
         \u_div/PartRem[19][16] , \u_div/PartRem[19][17] ,
         \u_div/PartRem[19][18] , \u_div/PartRem[19][19] ,
         \u_div/PartRem[19][20] , \u_div/PartRem[19][21] ,
         \u_div/PartRem[19][22] , \u_div/PartRem[19][23] ,
         \u_div/PartRem[19][24] , \u_div/PartRem[20][1] ,
         \u_div/PartRem[20][2] , \u_div/PartRem[20][3] ,
         \u_div/PartRem[20][4] , \u_div/PartRem[20][5] ,
         \u_div/PartRem[20][6] , \u_div/PartRem[20][7] ,
         \u_div/PartRem[20][8] , \u_div/PartRem[20][9] ,
         \u_div/PartRem[20][10] , \u_div/PartRem[20][11] ,
         \u_div/PartRem[20][12] , \u_div/PartRem[20][13] ,
         \u_div/PartRem[20][14] , \u_div/PartRem[20][15] ,
         \u_div/PartRem[20][16] , \u_div/PartRem[20][17] ,
         \u_div/PartRem[20][18] , \u_div/PartRem[20][19] ,
         \u_div/PartRem[20][20] , \u_div/PartRem[20][21] ,
         \u_div/PartRem[20][22] , \u_div/PartRem[20][24] ,
         \u_div/PartRem[21][1] , \u_div/PartRem[21][2] ,
         \u_div/PartRem[21][3] , \u_div/PartRem[21][4] ,
         \u_div/PartRem[21][5] , \u_div/PartRem[21][6] ,
         \u_div/PartRem[21][7] , \u_div/PartRem[21][8] ,
         \u_div/PartRem[21][9] , \u_div/PartRem[21][10] ,
         \u_div/PartRem[21][11] , \u_div/PartRem[21][12] ,
         \u_div/PartRem[21][13] , \u_div/PartRem[21][14] ,
         \u_div/PartRem[21][15] , \u_div/PartRem[21][16] ,
         \u_div/PartRem[21][17] , \u_div/PartRem[21][18] ,
         \u_div/PartRem[21][19] , \u_div/PartRem[21][20] ,
         \u_div/PartRem[21][21] , \u_div/PartRem[21][22] ,
         \u_div/PartRem[21][23] , \u_div/PartRem[21][24] ,
         \u_div/PartRem[22][1] , \u_div/PartRem[22][3] ,
         \u_div/PartRem[22][4] , \u_div/PartRem[22][5] ,
         \u_div/PartRem[22][6] , \u_div/PartRem[22][7] ,
         \u_div/PartRem[22][8] , \u_div/PartRem[22][9] ,
         \u_div/PartRem[22][10] , \u_div/PartRem[22][11] ,
         \u_div/PartRem[22][12] , \u_div/PartRem[22][13] ,
         \u_div/PartRem[22][14] , \u_div/PartRem[22][15] ,
         \u_div/PartRem[22][16] , \u_div/PartRem[22][17] ,
         \u_div/PartRem[22][18] , \u_div/PartRem[22][19] ,
         \u_div/PartRem[22][20] , \u_div/PartRem[22][21] ,
         \u_div/PartRem[22][22] , \u_div/PartRem[22][23] ,
         \u_div/PartRem[22][24] , \u_div/PartRem[23][2] ,
         \u_div/PartRem[23][3] , \u_div/PartRem[23][4] ,
         \u_div/PartRem[23][5] , \u_div/PartRem[23][6] ,
         \u_div/PartRem[23][7] , \u_div/PartRem[23][8] ,
         \u_div/PartRem[23][9] , \u_div/PartRem[23][10] ,
         \u_div/PartRem[23][11] , \u_div/PartRem[23][12] ,
         \u_div/PartRem[23][13] , \u_div/PartRem[23][14] ,
         \u_div/PartRem[23][15] , \u_div/PartRem[23][16] ,
         \u_div/PartRem[23][17] , \u_div/PartRem[23][18] ,
         \u_div/PartRem[23][19] , \u_div/PartRem[23][20] ,
         \u_div/PartRem[23][21] , \u_div/PartRem[23][22] ,
         \u_div/PartRem[23][23] , \u_div/PartRem[23][24] ,
         \u_div/PartRem[24][1] , \u_div/PartRem[24][2] ,
         \u_div/PartRem[24][3] , \u_div/PartRem[24][4] ,
         \u_div/PartRem[24][5] , \u_div/PartRem[24][6] ,
         \u_div/PartRem[24][7] , \u_div/PartRem[24][8] ,
         \u_div/PartRem[24][9] , \u_div/PartRem[24][10] ,
         \u_div/PartRem[24][11] , \u_div/PartRem[24][12] ,
         \u_div/PartRem[24][13] , \u_div/PartRem[24][14] ,
         \u_div/PartRem[24][15] , \u_div/PartRem[24][16] ,
         \u_div/PartRem[24][17] , \u_div/PartRem[24][18] ,
         \u_div/PartRem[24][19] , \u_div/PartRem[24][20] ,
         \u_div/PartRem[24][21] , \u_div/PartRem[24][22] ,
         \u_div/PartRem[24][23] , \u_div/PartRem[24][24] , \u_div/BInv[0] ,
         \u_div/BInv[3] , \u_div/BInv[4] , \u_div/BInv[5] , \u_div/BInv[6] ,
         \u_div/BInv[7] , \u_div/BInv[8] , \u_div/BInv[10] , \u_div/BInv[11] ,
         \u_div/BInv[12] , \u_div/BInv[13] , \u_div/BInv[14] ,
         \u_div/BInv[15] , \u_div/BInv[16] , \u_div/BInv[17] ,
         \u_div/BInv[18] , \u_div/BInv[19] , \u_div/BInv[20] ,
         \u_div/BInv[21] , \u_div/BInv[22] , n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n39, n40, n41, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n148, n150, n152, n154, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628;

  FADDX1_RVT \u_div/u_fa_PartRem_0_22_15  ( .A(\u_div/PartRem[23][15] ), .B(
        \u_div/BInv[15] ), .CI(\u_div/CryTmp[22][15] ), .CO(
        \u_div/CryTmp[22][16] ), .S(\u_div/SumTmp[22][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_20  ( .A(\u_div/PartRem[23][20] ), .B(
        \u_div/BInv[20] ), .CI(\u_div/CryTmp[22][20] ), .CO(
        \u_div/CryTmp[22][21] ), .S(\u_div/SumTmp[22][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_19  ( .A(\u_div/PartRem[22][19] ), .B(
        \u_div/BInv[19] ), .CI(\u_div/CryTmp[21][19] ), .CO(
        \u_div/CryTmp[21][20] ), .S(\u_div/SumTmp[21][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_17  ( .A(\u_div/PartRem[22][17] ), .B(
        \u_div/BInv[17] ), .CI(\u_div/CryTmp[21][17] ), .CO(
        \u_div/CryTmp[21][18] ), .S(\u_div/SumTmp[21][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_18  ( .A(\u_div/PartRem[22][18] ), .B(
        \u_div/BInv[18] ), .CI(\u_div/CryTmp[21][18] ), .CO(
        \u_div/CryTmp[21][19] ), .S(\u_div/SumTmp[21][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_16  ( .A(\u_div/PartRem[21][16] ), .B(
        \u_div/BInv[16] ), .CI(\u_div/CryTmp[20][16] ), .CO(
        \u_div/CryTmp[20][17] ), .S(\u_div/SumTmp[20][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_17  ( .A(\u_div/PartRem[21][17] ), .B(
        \u_div/BInv[17] ), .CI(\u_div/CryTmp[20][17] ), .CO(
        \u_div/CryTmp[20][18] ), .S(\u_div/SumTmp[20][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_17  ( .A(\u_div/PartRem[20][17] ), .B(
        \u_div/BInv[17] ), .CI(n35), .CO(\u_div/CryTmp[19][18] ), .S(
        \u_div/SumTmp[19][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_18  ( .A(\u_div/PartRem[19][18] ), .B(
        \u_div/BInv[18] ), .CI(\u_div/CryTmp[18][18] ), .CO(
        \u_div/CryTmp[18][19] ), .S(\u_div/SumTmp[18][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_19  ( .A(\u_div/PartRem[18][19] ), .B(
        \u_div/BInv[19] ), .CI(\u_div/CryTmp[17][19] ), .CO(
        \u_div/CryTmp[17][20] ), .S(\u_div/SumTmp[17][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_20  ( .A(\u_div/PartRem[17][20] ), .B(
        \u_div/BInv[20] ), .CI(\u_div/CryTmp[16][20] ), .CO(
        \u_div/CryTmp[16][21] ), .S(\u_div/SumTmp[16][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_21  ( .A(\u_div/PartRem[17][21] ), .B(
        \u_div/BInv[21] ), .CI(\u_div/CryTmp[16][21] ), .CO(
        \u_div/CryTmp[16][22] ), .S(\u_div/SumTmp[16][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_21  ( .A(\u_div/PartRem[16][21] ), .B(
        \u_div/BInv[21] ), .CI(\u_div/CryTmp[15][21] ), .CO(
        \u_div/CryTmp[15][22] ), .S(\u_div/SumTmp[15][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_22  ( .A(\u_div/PartRem[16][22] ), .B(
        \u_div/BInv[22] ), .CI(\u_div/CryTmp[15][22] ), .CO(
        \u_div/CryTmp[15][23] ), .S(\u_div/SumTmp[15][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_18  ( .A(\u_div/PartRem[18][18] ), .B(
        \u_div/BInv[18] ), .CI(\u_div/CryTmp[17][18] ), .CO(
        \u_div/CryTmp[17][19] ), .S(\u_div/SumTmp[17][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_16  ( .A(\u_div/PartRem[18][16] ), .B(
        \u_div/BInv[16] ), .CI(\u_div/CryTmp[17][16] ), .CO(
        \u_div/CryTmp[17][17] ), .S(\u_div/SumTmp[17][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_17  ( .A(\u_div/PartRem[18][17] ), .B(
        \u_div/BInv[17] ), .CI(\u_div/CryTmp[17][17] ), .CO(
        \u_div/CryTmp[17][18] ), .S(\u_div/SumTmp[17][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_3  ( .A(\u_div/PartRem[18][3] ), .B(
        \u_div/BInv[3] ), .CI(\u_div/CryTmp[17][3] ), .CO(
        \u_div/CryTmp[17][4] ), .S(\u_div/SumTmp[17][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_5  ( .A(\u_div/PartRem[17][5] ), .B(
        \u_div/BInv[5] ), .CI(\u_div/CryTmp[16][5] ), .CO(
        \u_div/CryTmp[16][6] ), .S(\u_div/SumTmp[16][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_4  ( .A(\u_div/PartRem[17][4] ), .B(
        \u_div/BInv[4] ), .CI(\u_div/CryTmp[16][4] ), .CO(
        \u_div/CryTmp[16][5] ), .S(\u_div/SumTmp[16][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_19  ( .A(\u_div/PartRem[16][19] ), .B(
        \u_div/BInv[19] ), .CI(\u_div/CryTmp[15][19] ), .CO(
        \u_div/CryTmp[15][20] ), .S(\u_div/SumTmp[15][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_17  ( .A(\u_div/PartRem[16][17] ), .B(
        \u_div/BInv[17] ), .CI(\u_div/CryTmp[15][17] ), .CO(
        \u_div/CryTmp[15][18] ), .S(\u_div/SumTmp[15][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_18  ( .A(\u_div/PartRem[16][18] ), .B(
        \u_div/BInv[18] ), .CI(n84), .CO(\u_div/CryTmp[15][19] ), .S(
        \u_div/SumTmp[15][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_5  ( .A(\u_div/PartRem[16][5] ), .B(
        \u_div/BInv[5] ), .CI(\u_div/CryTmp[15][5] ), .CO(
        \u_div/CryTmp[15][6] ), .S(\u_div/SumTmp[15][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_8  ( .A(\u_div/PartRem[15][8] ), .B(
        \u_div/BInv[8] ), .CI(\u_div/CryTmp[14][8] ), .CO(
        \u_div/CryTmp[14][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_6  ( .A(\u_div/PartRem[15][6] ), .B(
        \u_div/BInv[6] ), .CI(\u_div/CryTmp[14][6] ), .CO(
        \u_div/CryTmp[14][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_7  ( .A(\u_div/PartRem[15][7] ), .B(
        \u_div/BInv[7] ), .CI(\u_div/CryTmp[14][7] ), .CO(
        \u_div/CryTmp[14][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_16  ( .A(\u_div/PartRem[24][16] ), .B(
        \u_div/BInv[16] ), .CI(\u_div/CryTmp[23][16] ), .CO(
        \u_div/CryTmp[23][17] ), .S(\u_div/SumTmp[23][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_14  ( .A(\u_div/PartRem[24][14] ), .B(
        \u_div/BInv[14] ), .CI(\u_div/CryTmp[23][14] ), .CO(
        \u_div/CryTmp[23][15] ), .S(\u_div/SumTmp[23][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_15  ( .A(\u_div/PartRem[24][15] ), .B(
        \u_div/BInv[15] ), .CI(\u_div/CryTmp[23][15] ), .CO(
        \u_div/CryTmp[23][16] ), .S(\u_div/SumTmp[23][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_9  ( .A(a[33]), .B(n132), .CI(
        \u_div/CryTmp[24][9] ), .CO(\u_div/CryTmp[24][10] ), .S(
        \u_div/SumTmp[24][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_10  ( .A(a[34]), .B(\u_div/BInv[10] ), 
        .CI(\u_div/CryTmp[24][10] ), .CO(\u_div/CryTmp[24][11] ), .S(
        \u_div/SumTmp[24][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_14  ( .A(a[38]), .B(\u_div/BInv[14] ), 
        .CI(\u_div/CryTmp[24][14] ), .CO(\u_div/CryTmp[24][15] ), .S(
        \u_div/SumTmp[24][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_15  ( .A(a[39]), .B(\u_div/BInv[15] ), 
        .CI(\u_div/CryTmp[24][15] ), .CO(\u_div/CryTmp[24][16] ), .S(
        \u_div/SumTmp[24][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_18  ( .A(a[42]), .B(\u_div/BInv[18] ), 
        .CI(\u_div/CryTmp[24][18] ), .CO(\u_div/CryTmp[24][19] ), .S(
        \u_div/SumTmp[24][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_19  ( .A(a[43]), .B(\u_div/BInv[19] ), 
        .CI(\u_div/CryTmp[24][19] ), .CO(\u_div/CryTmp[24][20] ), .S(
        \u_div/SumTmp[24][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_1  ( .A(a[25]), .B(n139), .CI(
        \u_div/CryTmp[24][1] ), .CO(\u_div/CryTmp[24][2] ), .S(
        \u_div/SumTmp[24][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_17  ( .A(\u_div/PartRem[23][17] ), .B(
        \u_div/BInv[17] ), .CI(\u_div/CryTmp[22][17] ), .CO(
        \u_div/CryTmp[22][18] ), .S(\u_div/SumTmp[22][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_18  ( .A(\u_div/PartRem[23][18] ), .B(
        \u_div/BInv[18] ), .CI(\u_div/CryTmp[22][18] ), .CO(
        \u_div/CryTmp[22][19] ), .S(\u_div/SumTmp[22][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_21  ( .A(\u_div/PartRem[22][21] ), .B(
        n76), .CI(\u_div/BInv[21] ), .CO(\u_div/CryTmp[21][22] ), .S(
        \u_div/SumTmp[21][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_22  ( .A(\u_div/PartRem[22][22] ), .B(
        \u_div/BInv[22] ), .CI(\u_div/CryTmp[21][22] ), .CO(
        \u_div/CryTmp[21][23] ), .S(\u_div/SumTmp[21][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_16  ( .A(\u_div/PartRem[22][16] ), .B(
        \u_div/BInv[16] ), .CI(\u_div/CryTmp[21][16] ), .CO(
        \u_div/CryTmp[21][17] ), .S(\u_div/SumTmp[21][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_22  ( .A(\u_div/PartRem[21][22] ), .B(
        \u_div/BInv[22] ), .CI(n95), .CO(\u_div/CryTmp[20][23] ), .S(
        \u_div/SumTmp[20][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_20  ( .A(\u_div/PartRem[20][20] ), .B(
        \u_div/BInv[20] ), .CI(\u_div/CryTmp[19][20] ), .CO(
        \u_div/CryTmp[19][21] ), .S(\u_div/SumTmp[19][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_21  ( .A(\u_div/PartRem[20][21] ), .B(
        \u_div/BInv[21] ), .CI(\u_div/CryTmp[19][21] ), .CO(
        \u_div/CryTmp[19][22] ), .S(\u_div/SumTmp[19][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_22  ( .A(\u_div/PartRem[19][22] ), .B(
        \u_div/BInv[22] ), .CI(\u_div/CryTmp[18][22] ), .CO(
        \u_div/CryTmp[18][23] ), .S(\u_div/SumTmp[18][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_21  ( .A(\u_div/PartRem[18][21] ), .B(
        \u_div/BInv[21] ), .CI(n86), .CO(\u_div/CryTmp[17][22] ), .S(
        \u_div/SumTmp[17][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_22  ( .A(\u_div/PartRem[18][22] ), .B(
        \u_div/BInv[22] ), .CI(\u_div/CryTmp[17][22] ), .CO(
        \u_div/CryTmp[17][23] ), .S(\u_div/SumTmp[17][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_11  ( .A(\u_div/PartRem[18][11] ), .B(
        \u_div/BInv[11] ), .CI(\u_div/CryTmp[17][11] ), .CO(
        \u_div/CryTmp[17][12] ), .S(\u_div/SumTmp[17][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_12  ( .A(\u_div/PartRem[18][12] ), .B(
        \u_div/BInv[12] ), .CI(\u_div/CryTmp[17][12] ), .CO(
        \u_div/CryTmp[17][13] ), .S(\u_div/SumTmp[17][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_19  ( .A(\u_div/PartRem[17][19] ), .B(
        \u_div/BInv[19] ), .CI(n78), .CO(\u_div/CryTmp[16][20] ), .S(
        \u_div/SumTmp[16][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_8  ( .A(\u_div/PartRem[17][8] ), .B(
        \u_div/BInv[8] ), .CI(\u_div/CryTmp[16][8] ), .CO(
        \u_div/CryTmp[16][9] ), .S(\u_div/SumTmp[16][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_9  ( .A(\u_div/PartRem[17][9] ), .B(n132), .CI(\u_div/CryTmp[16][9] ), .CO(\u_div/CryTmp[16][10] ), .S(
        \u_div/SumTmp[16][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_20  ( .A(\u_div/PartRem[16][20] ), .B(
        \u_div/BInv[20] ), .CI(\u_div/CryTmp[15][20] ), .CO(
        \u_div/CryTmp[15][21] ), .S(\u_div/SumTmp[15][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_13  ( .A(\u_div/PartRem[16][13] ), .B(
        \u_div/BInv[13] ), .CI(n18), .CO(\u_div/CryTmp[15][14] ), .S(
        \u_div/SumTmp[15][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_6  ( .A(\u_div/PartRem[16][6] ), .B(
        \u_div/BInv[6] ), .CI(\u_div/CryTmp[15][6] ), .CO(
        \u_div/CryTmp[15][7] ), .S(\u_div/SumTmp[15][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_14  ( .A(\u_div/PartRem[15][14] ), .B(
        \u_div/BInv[14] ), .CI(\u_div/CryTmp[14][14] ), .CO(
        \u_div/CryTmp[14][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_15  ( .A(\u_div/PartRem[15][15] ), .B(
        \u_div/BInv[15] ), .CI(\u_div/CryTmp[14][15] ), .CO(
        \u_div/CryTmp[14][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_14  ( .A(\u_div/PartRem[16][14] ), .B(
        \u_div/BInv[14] ), .CI(\u_div/CryTmp[15][14] ), .CO(
        \u_div/CryTmp[15][15] ), .S(\u_div/SumTmp[15][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_15  ( .A(\u_div/PartRem[16][15] ), .B(
        \u_div/BInv[15] ), .CI(\u_div/CryTmp[15][15] ), .CO(
        \u_div/CryTmp[15][16] ), .S(\u_div/SumTmp[15][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_21  ( .A(\u_div/PartRem[24][21] ), .B(
        \u_div/BInv[21] ), .CI(n2), .CO(\u_div/CryTmp[23][22] ), .S(
        \u_div/SumTmp[23][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_22  ( .A(\u_div/PartRem[24][22] ), .B(
        \u_div/BInv[22] ), .CI(n33), .CO(\u_div/CryTmp[23][23] ), .S(
        \u_div/SumTmp[23][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_2  ( .A(a[26]), .B(n137), .CI(
        \u_div/CryTmp[24][2] ), .CO(\u_div/CryTmp[24][3] ), .S(
        \u_div/SumTmp[24][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_3  ( .A(a[27]), .B(n136), .CI(
        \u_div/CryTmp[24][3] ), .CO(\u_div/CryTmp[24][4] ), .S(
        \u_div/SumTmp[24][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_16  ( .A(\u_div/PartRem[23][16] ), .B(
        \u_div/BInv[16] ), .CI(\u_div/CryTmp[22][16] ), .CO(
        \u_div/CryTmp[22][17] ), .S(\u_div/SumTmp[22][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_19  ( .A(\u_div/PartRem[23][19] ), .B(
        \u_div/BInv[19] ), .CI(\u_div/CryTmp[22][19] ), .CO(
        \u_div/CryTmp[22][20] ), .S(\u_div/SumTmp[22][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_19  ( .A(\u_div/CryTmp[19][19] ), .B(
        \u_div/BInv[19] ), .CI(\u_div/PartRem[20][19] ), .CO(
        \u_div/CryTmp[19][20] ), .S(\u_div/SumTmp[19][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_20  ( .A(\u_div/PartRem[19][20] ), .B(
        \u_div/BInv[20] ), .CI(n8), .CO(\u_div/CryTmp[18][21] ), .S(
        \u_div/SumTmp[18][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_17  ( .A(\u_div/PartRem[19][17] ), .B(
        \u_div/BInv[17] ), .CI(n57), .CO(\u_div/CryTmp[18][18] ), .S(
        \u_div/SumTmp[18][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_9  ( .A(\u_div/PartRem[18][9] ), .B(n132), .CI(\u_div/CryTmp[17][9] ), .CO(\u_div/CryTmp[17][10] ), .S(
        \u_div/SumTmp[17][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_10  ( .A(\u_div/PartRem[18][10] ), .B(
        \u_div/BInv[10] ), .CI(\u_div/CryTmp[17][10] ), .CO(
        \u_div/CryTmp[17][11] ), .S(\u_div/SumTmp[17][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_5  ( .A(\u_div/PartRem[18][5] ), .B(
        \u_div/BInv[5] ), .CI(\u_div/CryTmp[17][5] ), .CO(
        \u_div/CryTmp[17][6] ), .S(\u_div/SumTmp[17][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_6  ( .A(\u_div/PartRem[18][6] ), .B(n133), .CI(\u_div/CryTmp[17][6] ), .CO(\u_div/CryTmp[17][7] ), .S(
        \u_div/SumTmp[17][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_17  ( .A(\u_div/PartRem[17][17] ), .B(
        n72), .CI(\u_div/BInv[17] ), .CO(\u_div/CryTmp[16][18] ), .S(
        \u_div/SumTmp[16][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_11  ( .A(\u_div/PartRem[17][11] ), .B(
        \u_div/BInv[11] ), .CI(\u_div/CryTmp[16][11] ), .CO(
        \u_div/CryTmp[16][12] ), .S(\u_div/SumTmp[16][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_12  ( .A(\u_div/PartRem[17][12] ), .B(
        \u_div/BInv[12] ), .CI(\u_div/CryTmp[16][12] ), .CO(
        \u_div/CryTmp[16][13] ), .S(\u_div/SumTmp[16][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_8  ( .A(\u_div/PartRem[16][8] ), .B(
        \u_div/BInv[8] ), .CI(\u_div/CryTmp[15][8] ), .CO(
        \u_div/CryTmp[15][9] ), .S(\u_div/SumTmp[15][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_9  ( .A(\u_div/PartRem[16][9] ), .B(n132), .CI(\u_div/CryTmp[15][9] ), .CO(\u_div/CryTmp[15][10] ), .S(
        \u_div/SumTmp[15][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_19  ( .A(\u_div/PartRem[15][19] ), .B(
        \u_div/BInv[19] ), .CI(n22), .CO(\u_div/CryTmp[14][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_20  ( .A(\u_div/PartRem[15][20] ), .B(
        \u_div/BInv[20] ), .CI(\u_div/CryTmp[14][20] ), .CO(
        \u_div/CryTmp[14][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_9  ( .A(\u_div/PartRem[15][9] ), .B(n132), .CI(\u_div/CryTmp[14][9] ), .CO(\u_div/CryTmp[14][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_10  ( .A(\u_div/PartRem[15][10] ), .B(
        \u_div/BInv[10] ), .CI(\u_div/CryTmp[14][10] ), .CO(
        \u_div/CryTmp[14][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_19  ( .A(\u_div/PartRem[24][19] ), .B(
        \u_div/BInv[19] ), .CI(\u_div/CryTmp[23][19] ), .CO(
        \u_div/CryTmp[23][20] ), .S(\u_div/SumTmp[23][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_20  ( .A(\u_div/PartRem[24][20] ), .B(
        \u_div/BInv[20] ), .CI(\u_div/CryTmp[23][20] ), .CO(
        \u_div/CryTmp[23][21] ), .S(\u_div/SumTmp[23][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_17  ( .A(\u_div/PartRem[24][17] ), .B(
        \u_div/BInv[17] ), .CI(\u_div/CryTmp[23][17] ), .CO(
        \u_div/CryTmp[23][18] ), .S(\u_div/SumTmp[23][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_12  ( .A(a[36]), .B(\u_div/BInv[12] ), 
        .CI(n12), .CO(\u_div/CryTmp[24][13] ), .S(\u_div/SumTmp[24][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_13  ( .A(a[37]), .B(\u_div/BInv[13] ), 
        .CI(\u_div/CryTmp[24][13] ), .CO(\u_div/CryTmp[24][14] ), .S(
        \u_div/SumTmp[24][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_7  ( .A(a[31]), .B(\u_div/BInv[7] ), 
        .CI(\u_div/CryTmp[24][7] ), .CO(\u_div/CryTmp[24][8] ), .S(
        \u_div/SumTmp[24][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_8  ( .A(a[32]), .B(\u_div/BInv[8] ), 
        .CI(\u_div/CryTmp[24][8] ), .CO(\u_div/CryTmp[24][9] ), .S(
        \u_div/SumTmp[24][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_22  ( .A(\u_div/PartRem[23][22] ), .B(
        \u_div/BInv[22] ), .CI(n91), .CO(\u_div/CryTmp[22][23] ), .S(
        \u_div/SumTmp[22][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_22  ( .A(\u_div/PartRem[20][22] ), .B(
        \u_div/BInv[22] ), .CI(\u_div/CryTmp[19][22] ), .CO(
        \u_div/CryTmp[19][23] ), .S(\u_div/SumTmp[19][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_7  ( .A(\u_div/PartRem[18][7] ), .B(
        \u_div/BInv[7] ), .CI(\u_div/CryTmp[17][7] ), .CO(
        \u_div/CryTmp[17][8] ), .S(\u_div/SumTmp[17][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_8  ( .A(\u_div/PartRem[18][8] ), .B(
        \u_div/BInv[8] ), .CI(\u_div/CryTmp[17][8] ), .CO(
        \u_div/CryTmp[17][9] ), .S(\u_div/SumTmp[17][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_10  ( .A(\u_div/PartRem[17][10] ), .B(
        \u_div/BInv[10] ), .CI(\u_div/CryTmp[16][10] ), .CO(
        \u_div/CryTmp[16][11] ), .S(\u_div/SumTmp[16][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_11  ( .A(\u_div/PartRem[16][11] ), .B(
        \u_div/BInv[11] ), .CI(\u_div/CryTmp[15][11] ), .CO(
        \u_div/CryTmp[15][12] ), .S(\u_div/SumTmp[15][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_12  ( .A(\u_div/PartRem[15][12] ), .B(
        \u_div/BInv[12] ), .CI(\u_div/CryTmp[14][12] ), .CO(
        \u_div/CryTmp[14][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_13  ( .A(\u_div/PartRem[15][13] ), .B(
        \u_div/BInv[13] ), .CI(\u_div/CryTmp[14][13] ), .CO(
        \u_div/CryTmp[14][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_6  ( .A(a[30]), .B(n133), .CI(
        \u_div/CryTmp[24][6] ), .CO(\u_div/CryTmp[24][7] ), .S(
        \u_div/SumTmp[24][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_4  ( .A(a[28]), .B(n135), .CI(
        \u_div/CryTmp[24][4] ), .CO(\u_div/CryTmp[24][5] ), .S(
        \u_div/SumTmp[24][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_5  ( .A(a[29]), .B(n134), .CI(
        \u_div/CryTmp[24][5] ), .CO(\u_div/CryTmp[24][6] ), .S(
        \u_div/SumTmp[24][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_18  ( .A(\u_div/PartRem[24][18] ), .B(
        \u_div/BInv[18] ), .CI(\u_div/CryTmp[23][18] ), .CO(
        \u_div/CryTmp[23][19] ), .S(\u_div/SumTmp[23][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_12  ( .A(\u_div/PartRem[24][12] ), .B(
        \u_div/BInv[12] ), .CI(n14), .CO(\u_div/CryTmp[23][13] ), .S(
        \u_div/SumTmp[23][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_11  ( .A(\u_div/PartRem[24][11] ), .B(
        \u_div/BInv[11] ), .CI(\u_div/CryTmp[23][11] ), .CO(
        \u_div/CryTmp[23][12] ), .S(\u_div/SumTmp[23][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_10  ( .A(\u_div/PartRem[24][10] ), .B(
        \u_div/BInv[10] ), .CI(\u_div/CryTmp[23][10] ), .CO(
        \u_div/CryTmp[23][11] ), .S(\u_div/SumTmp[23][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_13  ( .A(\u_div/PartRem[24][13] ), .B(
        \u_div/BInv[13] ), .CI(\u_div/CryTmp[23][13] ), .CO(
        \u_div/CryTmp[23][14] ), .S(\u_div/SumTmp[23][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_1  ( .A(\u_div/PartRem[24][1] ), .B(n139), .CI(\u_div/CryTmp[23][1] ), .CO(\u_div/CryTmp[23][2] ), .S(
        \u_div/SumTmp[23][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_21  ( .A(a[45]), .B(\u_div/BInv[21] ), 
        .CI(n80), .CO(\u_div/CryTmp[24][22] ), .S(\u_div/SumTmp[24][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_17  ( .A(a[41]), .B(\u_div/BInv[17] ), 
        .CI(n16), .CO(\u_div/CryTmp[24][18] ), .S(\u_div/SumTmp[24][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_10  ( .A(\u_div/PartRem[16][10] ), .B(
        \u_div/BInv[10] ), .CI(\u_div/CryTmp[15][10] ), .CO(
        \u_div/CryTmp[15][11] ), .S(\u_div/SumTmp[15][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_15  ( .A(\u_div/PartRem[19][15] ), .B(
        \u_div/BInv[15] ), .CI(\u_div/CryTmp[18][15] ), .CO(
        \u_div/CryTmp[18][16] ), .S(\u_div/SumTmp[18][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_18  ( .A(\u_div/PartRem[21][18] ), .B(
        \u_div/BInv[18] ), .CI(\u_div/CryTmp[20][18] ), .CO(
        \u_div/CryTmp[20][19] ), .S(\u_div/SumTmp[20][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_19  ( .A(\u_div/PartRem[21][19] ), .B(
        \u_div/BInv[19] ), .CI(\u_div/CryTmp[20][19] ), .CO(
        \u_div/CryTmp[20][20] ), .S(\u_div/SumTmp[20][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_15  ( .A(\u_div/PartRem[22][15] ), .B(
        \u_div/BInv[15] ), .CI(\u_div/CryTmp[21][15] ), .CO(
        \u_div/CryTmp[21][16] ), .S(\u_div/SumTmp[21][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_11  ( .A(\u_div/PartRem[15][11] ), .B(
        \u_div/BInv[11] ), .CI(\u_div/CryTmp[14][11] ), .CO(
        \u_div/CryTmp[14][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_13  ( .A(\u_div/PartRem[20][13] ), .B(
        \u_div/BInv[13] ), .CI(\u_div/CryTmp[19][13] ), .CO(
        \u_div/CryTmp[19][14] ), .S(\u_div/SumTmp[19][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_12  ( .A(\u_div/PartRem[20][12] ), .B(
        \u_div/BInv[12] ), .CI(\u_div/CryTmp[19][12] ), .CO(
        \u_div/CryTmp[19][13] ), .S(\u_div/SumTmp[19][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_11  ( .A(\u_div/PartRem[20][11] ), .B(
        \u_div/BInv[11] ), .CI(\u_div/CryTmp[19][11] ), .CO(
        \u_div/CryTmp[19][12] ), .S(\u_div/SumTmp[19][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_14  ( .A(\u_div/PartRem[20][14] ), .B(
        \u_div/BInv[14] ), .CI(\u_div/CryTmp[19][14] ), .CO(
        \u_div/CryTmp[19][15] ), .S(\u_div/SumTmp[19][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_15  ( .A(\u_div/PartRem[20][15] ), .B(
        \u_div/BInv[15] ), .CI(\u_div/CryTmp[19][15] ), .CO(
        \u_div/CryTmp[19][16] ), .S(\u_div/SumTmp[19][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_10  ( .A(\u_div/PartRem[19][10] ), .B(
        \u_div/BInv[10] ), .CI(\u_div/CryTmp[18][10] ), .CO(
        \u_div/CryTmp[18][11] ), .S(\u_div/SumTmp[18][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_14  ( .A(\u_div/PartRem[19][14] ), .B(
        \u_div/BInv[14] ), .CI(n6), .CO(\u_div/CryTmp[18][15] ), .S(
        \u_div/SumTmp[18][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_13  ( .A(\u_div/PartRem[19][13] ), .B(
        \u_div/BInv[13] ), .CI(n74), .CO(\u_div/CryTmp[18][14] ), .S(
        \u_div/SumTmp[18][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_13  ( .A(\u_div/PartRem[17][13] ), .B(
        \u_div/BInv[13] ), .CI(\u_div/CryTmp[16][13] ), .CO(
        \u_div/CryTmp[16][14] ), .S(\u_div/SumTmp[16][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_17  ( .A(\u_div/PartRem[15][17] ), .B(
        \u_div/BInv[17] ), .CI(\u_div/CryTmp[14][17] ), .CO(
        \u_div/CryTmp[14][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_14  ( .A(\u_div/PartRem[18][14] ), .B(
        \u_div/BInv[14] ), .CI(\u_div/CryTmp[17][14] ), .CO(
        \u_div/CryTmp[17][15] ), .S(\u_div/SumTmp[17][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_13  ( .A(\u_div/PartRem[18][13] ), .B(
        \u_div/BInv[13] ), .CI(\u_div/CryTmp[17][13] ), .CO(
        \u_div/CryTmp[17][14] ), .S(\u_div/SumTmp[17][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_15  ( .A(\u_div/PartRem[18][15] ), .B(
        \u_div/BInv[15] ), .CI(n10), .CO(\u_div/CryTmp[17][16] ), .S(
        \u_div/SumTmp[17][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_14  ( .A(\u_div/PartRem[17][14] ), .B(
        \u_div/BInv[14] ), .CI(\u_div/CryTmp[16][14] ), .CO(
        \u_div/CryTmp[16][15] ), .S(\u_div/SumTmp[16][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_15  ( .A(\u_div/PartRem[17][15] ), .B(
        \u_div/BInv[15] ), .CI(\u_div/CryTmp[16][15] ), .CO(
        \u_div/CryTmp[16][16] ), .S(\u_div/SumTmp[16][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_10  ( .A(\u_div/PartRem[21][10] ), .B(
        \u_div/BInv[10] ), .CI(\u_div/CryTmp[20][10] ), .CO(
        \u_div/CryTmp[20][11] ), .S(\u_div/SumTmp[20][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_11  ( .A(\u_div/PartRem[21][11] ), .B(
        \u_div/BInv[11] ), .CI(\u_div/CryTmp[20][11] ), .CO(
        \u_div/CryTmp[20][12] ), .S(\u_div/SumTmp[20][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_13  ( .A(\u_div/PartRem[21][13] ), .B(
        \u_div/BInv[13] ), .CI(n45), .CO(\u_div/CryTmp[20][14] ), .S(
        \u_div/SumTmp[20][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_14  ( .A(\u_div/PartRem[21][14] ), .B(
        \u_div/BInv[14] ), .CI(\u_div/CryTmp[20][14] ), .CO(
        \u_div/CryTmp[20][15] ), .S(\u_div/SumTmp[20][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_10  ( .A(\u_div/PartRem[22][10] ), .B(
        \u_div/BInv[10] ), .CI(\u_div/CryTmp[21][10] ), .CO(
        \u_div/CryTmp[21][11] ), .S(\u_div/SumTmp[21][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_12  ( .A(\u_div/PartRem[22][12] ), .B(
        \u_div/BInv[12] ), .CI(n4), .CO(\u_div/CryTmp[21][13] ), .S(
        \u_div/SumTmp[21][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_13  ( .A(\u_div/PartRem[22][13] ), .B(
        \u_div/BInv[13] ), .CI(\u_div/CryTmp[21][13] ), .CO(
        \u_div/CryTmp[21][14] ), .S(\u_div/SumTmp[21][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_14  ( .A(\u_div/PartRem[22][14] ), .B(
        \u_div/BInv[14] ), .CI(\u_div/CryTmp[21][14] ), .CO(
        \u_div/CryTmp[21][15] ), .S(\u_div/SumTmp[21][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_10  ( .A(\u_div/PartRem[23][10] ), .B(
        \u_div/BInv[10] ), .CI(\u_div/CryTmp[22][10] ), .CO(
        \u_div/CryTmp[22][11] ), .S(\u_div/SumTmp[22][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_11  ( .A(\u_div/PartRem[23][11] ), .B(
        \u_div/BInv[11] ), .CI(\u_div/CryTmp[22][11] ), .CO(
        \u_div/CryTmp[22][12] ), .S(\u_div/SumTmp[22][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_13  ( .A(\u_div/PartRem[23][13] ), .B(
        \u_div/BInv[13] ), .CI(n89), .CO(\u_div/CryTmp[22][14] ), .S(
        \u_div/SumTmp[22][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_14  ( .A(\u_div/PartRem[23][14] ), .B(
        \u_div/BInv[14] ), .CI(\u_div/CryTmp[22][14] ), .CO(
        \u_div/CryTmp[22][15] ), .S(\u_div/SumTmp[22][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_9  ( .A(\u_div/PartRem[24][9] ), .B(n132), .CI(\u_div/CryTmp[23][9] ), .CO(\u_div/CryTmp[23][10] ), .S(
        \u_div/SumTmp[23][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_8  ( .A(\u_div/PartRem[24][8] ), .B(
        \u_div/BInv[8] ), .CI(\u_div/CryTmp[23][8] ), .CO(
        \u_div/CryTmp[23][9] ), .S(\u_div/SumTmp[23][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_7  ( .A(\u_div/PartRem[24][7] ), .B(
        \u_div/BInv[7] ), .CI(\u_div/CryTmp[23][7] ), .CO(
        \u_div/CryTmp[23][8] ), .S(\u_div/SumTmp[23][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_6  ( .A(\u_div/PartRem[24][6] ), .B(n133), .CI(\u_div/CryTmp[23][6] ), .CO(\u_div/CryTmp[23][7] ), .S(
        \u_div/SumTmp[23][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_5  ( .A(\u_div/PartRem[24][5] ), .B(n134), .CI(\u_div/CryTmp[23][5] ), .CO(\u_div/CryTmp[23][6] ), .S(
        \u_div/SumTmp[23][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_4  ( .A(\u_div/PartRem[24][4] ), .B(n135), .CI(\u_div/CryTmp[23][4] ), .CO(\u_div/CryTmp[23][5] ), .S(
        \u_div/SumTmp[23][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_3  ( .A(\u_div/PartRem[24][3] ), .B(n136), .CI(\u_div/CryTmp[23][3] ), .CO(\u_div/CryTmp[23][4] ), .S(
        \u_div/SumTmp[23][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_2  ( .A(\u_div/PartRem[24][2] ), .B(n137), .CI(\u_div/CryTmp[23][2] ), .CO(\u_div/CryTmp[23][3] ), .S(
        \u_div/SumTmp[23][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_1  ( .A(n140), .B(n51), .CI(
        \u_div/CryTmp[23][1] ), .CO(\u_div/CryTmp[20][2] ), .S(
        \u_div/SumTmp[20][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_1  ( .A(\u_div/PartRem[22][1] ), .B(n140), .CI(\u_div/CryTmp[23][1] ), .CO(\u_div/CryTmp[21][2] ), .S(
        \u_div/SumTmp[21][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_2  ( .A(\u_div/PartRem[21][2] ), .B(n138), .CI(\u_div/CryTmp[20][2] ), .CO(\u_div/CryTmp[20][3] ), .S(
        \u_div/SumTmp[20][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_2  ( .A(n55), .B(n138), .CI(
        \u_div/CryTmp[19][2] ), .CO(\u_div/CryTmp[19][3] ), .S(
        \u_div/SumTmp[19][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_3  ( .A(\u_div/PartRem[20][3] ), .B(
        \u_div/BInv[3] ), .CI(\u_div/CryTmp[19][3] ), .CO(
        \u_div/CryTmp[19][4] ), .S(\u_div/SumTmp[19][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_1  ( .A(n60), .B(n140), .CI(
        \u_div/CryTmp[23][1] ), .CO(\u_div/CryTmp[19][2] ), .S(
        \u_div/SumTmp[19][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_3  ( .A(\u_div/PartRem[19][3] ), .B(
        \u_div/BInv[3] ), .CI(\u_div/CryTmp[18][3] ), .CO(
        \u_div/CryTmp[18][4] ), .S(\u_div/SumTmp[18][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_2  ( .A(\u_div/PartRem[19][2] ), .B(n138), .CI(\u_div/CryTmp[18][2] ), .CO(\u_div/CryTmp[18][3] ), .S(
        \u_div/SumTmp[18][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_4  ( .A(\u_div/PartRem[19][4] ), .B(
        \u_div/BInv[4] ), .CI(\u_div/CryTmp[18][4] ), .CO(
        \u_div/CryTmp[18][5] ), .S(\u_div/SumTmp[18][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_1  ( .A(\u_div/PartRem[19][1] ), .B(n140), .CI(\u_div/CryTmp[23][1] ), .CO(\u_div/CryTmp[18][2] ), .S(
        \u_div/SumTmp[18][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_7  ( .A(\u_div/PartRem[17][7] ), .B(
        \u_div/BInv[7] ), .CI(\u_div/CryTmp[16][7] ), .CO(
        \u_div/CryTmp[16][8] ), .S(\u_div/SumTmp[16][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_7  ( .A(\u_div/PartRem[16][7] ), .B(
        \u_div/BInv[7] ), .CI(\u_div/CryTmp[15][7] ), .CO(
        \u_div/CryTmp[15][8] ), .S(\u_div/SumTmp[15][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_6  ( .A(\u_div/PartRem[17][6] ), .B(
        \u_div/BInv[6] ), .CI(\u_div/CryTmp[16][6] ), .CO(
        \u_div/CryTmp[16][7] ), .S(\u_div/SumTmp[16][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_4  ( .A(\u_div/PartRem[18][4] ), .B(
        \u_div/BInv[4] ), .CI(\u_div/CryTmp[17][4] ), .CO(
        \u_div/CryTmp[17][5] ), .S(\u_div/SumTmp[17][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_5  ( .A(\u_div/PartRem[15][5] ), .B(
        \u_div/BInv[5] ), .CI(\u_div/CryTmp[14][5] ), .CO(
        \u_div/CryTmp[14][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_2  ( .A(\u_div/PartRem[16][2] ), .B(n138), .CI(\u_div/CryTmp[15][2] ), .CO(\u_div/CryTmp[15][3] ), .S(
        \u_div/SumTmp[15][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_1  ( .A(n49), .B(n140), .CI(
        \u_div/CryTmp[23][1] ), .CO(\u_div/CryTmp[16][2] ), .S(
        \u_div/SumTmp[16][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_7  ( .A(\u_div/PartRem[20][7] ), .B(
        \u_div/BInv[7] ), .CI(\u_div/CryTmp[19][7] ), .CO(
        \u_div/CryTmp[19][8] ), .S(\u_div/SumTmp[19][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_8  ( .A(\u_div/PartRem[20][8] ), .B(
        \u_div/BInv[8] ), .CI(\u_div/CryTmp[19][8] ), .CO(
        \u_div/CryTmp[19][9] ), .S(\u_div/SumTmp[19][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_9  ( .A(\u_div/PartRem[20][9] ), .B(n132), .CI(\u_div/CryTmp[19][9] ), .CO(\u_div/CryTmp[19][10] ), .S(
        \u_div/SumTmp[19][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_6  ( .A(\u_div/PartRem[20][6] ), .B(
        \u_div/CryTmp[19][6] ), .CI(n133), .CO(\u_div/CryTmp[19][7] ), .S(
        \u_div/SumTmp[19][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_3  ( .A(\u_div/PartRem[16][3] ), .B(
        \u_div/BInv[3] ), .CI(\u_div/CryTmp[15][3] ), .CO(
        \u_div/CryTmp[15][4] ), .S(\u_div/SumTmp[15][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_4  ( .A(\u_div/PartRem[16][4] ), .B(
        \u_div/BInv[4] ), .CI(\u_div/CryTmp[15][4] ), .CO(
        \u_div/CryTmp[15][5] ), .S(\u_div/SumTmp[15][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_8  ( .A(\u_div/PartRem[19][8] ), .B(
        \u_div/BInv[8] ), .CI(\u_div/CryTmp[18][8] ), .CO(
        \u_div/CryTmp[18][9] ), .S(\u_div/SumTmp[18][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_7  ( .A(\u_div/PartRem[19][7] ), .B(
        \u_div/BInv[7] ), .CI(\u_div/CryTmp[18][7] ), .CO(
        \u_div/CryTmp[18][8] ), .S(\u_div/SumTmp[18][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_3  ( .A(\u_div/PartRem[15][3] ), .B(
        \u_div/BInv[3] ), .CI(\u_div/CryTmp[14][3] ), .CO(
        \u_div/CryTmp[14][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_4  ( .A(\u_div/PartRem[15][4] ), .B(
        \u_div/BInv[4] ), .CI(\u_div/CryTmp[14][4] ), .CO(
        \u_div/CryTmp[14][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_1  ( .A(n39), .B(n140), .CI(
        \u_div/CryTmp[23][1] ), .CO(\u_div/CryTmp[14][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_2  ( .A(\u_div/PartRem[15][2] ), .B(n138), .CI(\u_div/CryTmp[14][2] ), .CO(\u_div/CryTmp[14][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_6  ( .A(\u_div/PartRem[19][6] ), .B(n133), .CI(\u_div/CryTmp[18][6] ), .CO(\u_div/CryTmp[18][7] ), .S(
        \u_div/SumTmp[18][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_1  ( .A(\u_div/PartRem[18][1] ), .B(n140), .CI(\u_div/CryTmp[23][1] ), .CO(\u_div/CryTmp[17][2] ), .S(
        \u_div/SumTmp[17][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_2  ( .A(\u_div/PartRem[18][2] ), .B(n138), .CI(\u_div/CryTmp[17][2] ), .CO(\u_div/CryTmp[17][3] ), .S(
        \u_div/SumTmp[17][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_5  ( .A(\u_div/PartRem[20][5] ), .B(n134), .CI(\u_div/CryTmp[19][5] ), .CO(\u_div/CryTmp[19][6] ), .S(
        \u_div/SumTmp[19][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_2  ( .A(\u_div/PartRem[17][2] ), .B(n138), .CI(\u_div/CryTmp[16][2] ), .CO(\u_div/CryTmp[16][3] ), .S(
        \u_div/SumTmp[16][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_3  ( .A(\u_div/PartRem[17][3] ), .B(
        \u_div/BInv[3] ), .CI(\u_div/CryTmp[16][3] ), .CO(
        \u_div/CryTmp[16][4] ), .S(\u_div/SumTmp[16][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_6  ( .A(\u_div/PartRem[21][6] ), .B(n133), .CI(\u_div/CryTmp[20][6] ), .CO(\u_div/CryTmp[20][7] ), .S(
        \u_div/SumTmp[20][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_7  ( .A(\u_div/PartRem[21][7] ), .B(
        \u_div/BInv[7] ), .CI(\u_div/CryTmp[20][7] ), .CO(
        \u_div/CryTmp[20][8] ), .S(\u_div/SumTmp[20][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_8  ( .A(\u_div/PartRem[21][8] ), .B(
        \u_div/BInv[8] ), .CI(\u_div/CryTmp[20][8] ), .CO(
        \u_div/CryTmp[20][9] ), .S(\u_div/SumTmp[20][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_9  ( .A(\u_div/PartRem[21][9] ), .B(n132), .CI(\u_div/CryTmp[20][9] ), .CO(\u_div/CryTmp[20][10] ), .S(
        \u_div/SumTmp[20][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_4  ( .A(\u_div/PartRem[21][4] ), .B(n135), .CI(\u_div/CryTmp[20][4] ), .CO(\u_div/CryTmp[20][5] ), .S(
        \u_div/SumTmp[20][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_3  ( .A(\u_div/PartRem[22][3] ), .B(n136), .CI(\u_div/CryTmp[21][3] ), .CO(\u_div/CryTmp[21][4] ), .S(
        \u_div/SumTmp[21][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_4  ( .A(\u_div/PartRem[22][4] ), .B(n135), .CI(\u_div/CryTmp[21][4] ), .CO(\u_div/CryTmp[21][5] ), .S(
        \u_div/SumTmp[21][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_5  ( .A(\u_div/PartRem[22][5] ), .B(n134), .CI(\u_div/CryTmp[21][5] ), .CO(\u_div/CryTmp[21][6] ), .S(
        \u_div/SumTmp[21][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_6  ( .A(\u_div/PartRem[22][6] ), .B(n133), .CI(\u_div/CryTmp[21][6] ), .CO(\u_div/CryTmp[21][7] ), .S(
        \u_div/SumTmp[21][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_7  ( .A(\u_div/PartRem[22][7] ), .B(
        \u_div/BInv[7] ), .CI(\u_div/CryTmp[21][7] ), .CO(
        \u_div/CryTmp[21][8] ), .S(\u_div/SumTmp[21][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_8  ( .A(\u_div/PartRem[22][8] ), .B(
        \u_div/BInv[8] ), .CI(\u_div/CryTmp[21][8] ), .CO(
        \u_div/CryTmp[21][9] ), .S(\u_div/SumTmp[21][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_9  ( .A(\u_div/PartRem[22][9] ), .B(n132), .CI(\u_div/CryTmp[21][9] ), .CO(\u_div/CryTmp[21][10] ), .S(
        \u_div/SumTmp[21][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_2  ( .A(\u_div/PartRem[23][2] ), .B(n137), .CI(\u_div/CryTmp[22][2] ), .CO(\u_div/CryTmp[22][3] ), .S(
        \u_div/SumTmp[22][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_3  ( .A(\u_div/PartRem[23][3] ), .B(n136), .CI(\u_div/CryTmp[22][3] ), .CO(\u_div/CryTmp[22][4] ), .S(
        \u_div/SumTmp[22][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_4  ( .A(\u_div/PartRem[23][4] ), .B(n135), .CI(\u_div/CryTmp[22][4] ), .CO(\u_div/CryTmp[22][5] ), .S(
        \u_div/SumTmp[22][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_5  ( .A(\u_div/PartRem[23][5] ), .B(n134), .CI(\u_div/CryTmp[22][5] ), .CO(\u_div/CryTmp[22][6] ), .S(
        \u_div/SumTmp[22][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_6  ( .A(\u_div/PartRem[23][6] ), .B(n133), .CI(\u_div/CryTmp[22][6] ), .CO(\u_div/CryTmp[22][7] ), .S(
        \u_div/SumTmp[22][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_7  ( .A(\u_div/PartRem[23][7] ), .B(
        \u_div/BInv[7] ), .CI(\u_div/CryTmp[22][7] ), .CO(
        \u_div/CryTmp[22][8] ), .S(\u_div/SumTmp[22][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_8  ( .A(\u_div/PartRem[23][8] ), .B(
        \u_div/BInv[8] ), .CI(\u_div/CryTmp[22][8] ), .CO(
        \u_div/CryTmp[22][9] ), .S(\u_div/SumTmp[22][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_9  ( .A(\u_div/PartRem[23][9] ), .B(n132), .CI(\u_div/CryTmp[22][9] ), .CO(\u_div/CryTmp[22][10] ), .S(
        \u_div/SumTmp[22][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_5  ( .A(\u_div/PartRem[19][5] ), .B(n134), .CI(\u_div/CryTmp[18][5] ), .CO(\u_div/CryTmp[18][6] ), .S(
        \u_div/SumTmp[18][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_1  ( .A(\u_div/PartRem[16][1] ), .B(n140), .CI(\u_div/CryTmp[23][1] ), .CO(\u_div/CryTmp[15][2] ), .S(
        \u_div/SumTmp[15][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_4  ( .A(\u_div/PartRem[20][4] ), .B(n135), .CI(\u_div/CryTmp[19][4] ), .CO(\u_div/CryTmp[19][5] ), .S(
        \u_div/SumTmp[19][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_3  ( .A(\u_div/PartRem[21][3] ), .B(n136), .CI(\u_div/CryTmp[20][3] ), .CO(\u_div/CryTmp[20][4] ), .S(
        \u_div/SumTmp[20][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_2  ( .A(\u_div/CryTmp[21][2] ), .B(n138), 
        .CI(n52), .CO(\u_div/CryTmp[21][3] ), .S(\u_div/SumTmp[21][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_1  ( .A(n40), .B(n140), .CI(
        \u_div/CryTmp[23][1] ), .CO(\u_div/CryTmp[22][2] ), .S(
        \u_div/SumTmp[22][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_5  ( .A(\u_div/PartRem[21][5] ), .B(n134), .CI(\u_div/CryTmp[20][5] ), .CO(\u_div/CryTmp[20][6] ), .S(
        \u_div/SumTmp[20][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_16  ( .A(\u_div/PartRem[16][16] ), .B(
        \u_div/BInv[16] ), .CI(\u_div/CryTmp[15][16] ), .CO(
        \u_div/CryTmp[15][17] ), .S(\u_div/SumTmp[15][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_16  ( .A(\u_div/PartRem[15][16] ), .B(
        \u_div/BInv[16] ), .CI(\u_div/CryTmp[14][16] ), .CO(
        \u_div/CryTmp[14][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_21  ( .A(\u_div/PartRem[19][21] ), .B(
        \u_div/BInv[21] ), .CI(\u_div/CryTmp[18][21] ), .CO(
        \u_div/CryTmp[18][22] ), .S(\u_div/SumTmp[18][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_22  ( .A(\u_div/PartRem[15][22] ), .B(
        n93), .CI(\u_div/BInv[22] ), .CO(\u_div/CryTmp[14][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_22  ( .A(\u_div/PartRem[17][22] ), .B(
        \u_div/BInv[22] ), .CI(\u_div/CryTmp[16][22] ), .CO(
        \u_div/CryTmp[16][23] ), .S(\u_div/SumTmp[16][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_22  ( .A(a[46]), .B(\u_div/BInv[22] ), 
        .CI(n70), .CO(\u_div/CryTmp[24][24] ), .S(\u_div/SumTmp[24][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_20  ( .A(a[44]), .B(\u_div/BInv[20] ), 
        .CI(\u_div/CryTmp[24][20] ), .CO(\u_div/CryTmp[24][21] ), .S(
        \u_div/SumTmp[24][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_9  ( .A(\u_div/PartRem[19][9] ), .B(n132), .CI(\u_div/CryTmp[18][9] ), .CO(\u_div/CryTmp[18][10] ), .S(
        \u_div/SumTmp[18][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_18  ( .A(\u_div/PartRem[20][18] ), .B(
        \u_div/BInv[18] ), .CI(\u_div/CryTmp[19][18] ), .CO(
        \u_div/CryTmp[19][19] ), .S(\u_div/SumTmp[19][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_16  ( .A(\u_div/PartRem[19][16] ), .B(
        \u_div/BInv[16] ), .CI(\u_div/CryTmp[18][16] ), .CO(
        \u_div/CryTmp[18][17] ), .S(\u_div/SumTmp[18][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_15  ( .A(\u_div/PartRem[21][15] ), .B(
        \u_div/BInv[15] ), .CI(\u_div/CryTmp[20][15] ), .CO(
        \u_div/CryTmp[20][16] ), .S(\u_div/SumTmp[20][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_12  ( .A(\u_div/PartRem[23][12] ), .B(
        \u_div/BInv[12] ), .CI(\u_div/CryTmp[22][12] ), .CO(
        \u_div/CryTmp[22][13] ), .S(\u_div/SumTmp[22][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_21  ( .A(\u_div/PartRem[23][21] ), .B(
        \u_div/BInv[21] ), .CI(\u_div/CryTmp[22][21] ), .CO(
        \u_div/CryTmp[22][22] ), .S(\u_div/SumTmp[22][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_20  ( .A(\u_div/PartRem[21][20] ), .B(
        \u_div/BInv[20] ), .CI(\u_div/CryTmp[20][20] ), .CO(
        \u_div/CryTmp[20][21] ), .S(\u_div/SumTmp[20][20] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_18_12  ( .A(\u_div/PartRem[19][12] ), .B(
        \u_div/BInv[12] ), .CI(n20), .CO(\u_div/CryTmp[18][13] ), .S(
        \u_div/SumTmp[18][12] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_16_16  ( .A(\u_div/PartRem[17][16] ), .B(
        \u_div/BInv[16] ), .CI(\u_div/CryTmp[16][16] ), .CO(
        \u_div/CryTmp[16][17] ), .S(\u_div/SumTmp[16][16] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_14_18  ( .A(\u_div/PartRem[15][18] ), .B(
        \u_div/BInv[18] ), .CI(\u_div/CryTmp[14][18] ), .CO(
        \u_div/CryTmp[14][19] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_14_21  ( .A(\u_div/PartRem[15][21] ), .B(
        \u_div/BInv[21] ), .CI(\u_div/CryTmp[14][21] ), .CO(
        \u_div/CryTmp[14][22] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_21_20  ( .A(\u_div/PartRem[22][20] ), .B(
        \u_div/BInv[20] ), .CI(\u_div/CryTmp[21][20] ), .CO(
        \u_div/CryTmp[21][21] ), .S(\u_div/SumTmp[21][20] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_18_11  ( .A(\u_div/PartRem[19][11] ), .B(
        \u_div/BInv[11] ), .CI(\u_div/CryTmp[18][11] ), .CO(
        \u_div/CryTmp[18][12] ), .S(\u_div/SumTmp[18][11] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_17_20  ( .A(\u_div/PartRem[18][20] ), .B(
        \u_div/BInv[20] ), .CI(\u_div/CryTmp[17][20] ), .CO(
        \u_div/CryTmp[17][21] ), .S(\u_div/SumTmp[17][20] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_15_12  ( .A(\u_div/PartRem[16][12] ), .B(
        \u_div/BInv[12] ), .CI(\u_div/CryTmp[15][12] ), .CO(
        \u_div/CryTmp[15][13] ), .S(\u_div/SumTmp[15][12] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_24_16  ( .A(a[40]), .B(\u_div/BInv[16] ), 
        .CI(\u_div/CryTmp[24][16] ), .CO(\u_div/CryTmp[24][17] ), .S(
        \u_div/SumTmp[24][16] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_24_11  ( .A(a[35]), .B(\u_div/BInv[11] ), 
        .CI(\u_div/CryTmp[24][11] ), .CO(\u_div/CryTmp[24][12] ), .S(
        \u_div/SumTmp[24][11] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_19_16  ( .A(\u_div/PartRem[20][16] ), .B(
        \u_div/BInv[16] ), .CI(\u_div/CryTmp[19][16] ), .CO(
        \u_div/CryTmp[19][17] ), .S(\u_div/SumTmp[19][16] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_20_12  ( .A(\u_div/PartRem[21][12] ), .B(
        \u_div/BInv[12] ), .CI(\u_div/CryTmp[20][12] ), .CO(
        \u_div/CryTmp[20][13] ), .S(\u_div/SumTmp[20][12] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_18_19  ( .A(\u_div/PartRem[19][19] ), .B(
        \u_div/BInv[19] ), .CI(\u_div/CryTmp[18][19] ), .CO(
        \u_div/CryTmp[18][20] ), .S(\u_div/SumTmp[18][19] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_20_21  ( .A(\u_div/PartRem[21][21] ), .B(
        \u_div/BInv[21] ), .CI(\u_div/CryTmp[20][21] ), .CO(
        \u_div/CryTmp[20][22] ), .S(\u_div/SumTmp[20][21] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_21_11  ( .A(\u_div/PartRem[22][11] ), .B(
        \u_div/BInv[11] ), .CI(\u_div/CryTmp[21][11] ), .CO(
        \u_div/CryTmp[21][12] ), .S(\u_div/SumTmp[21][11] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_16_18  ( .A(\u_div/PartRem[17][18] ), .B(
        \u_div/BInv[18] ), .CI(\u_div/CryTmp[16][18] ), .CO(
        \u_div/CryTmp[16][19] ), .S(\u_div/SumTmp[16][18] ) );
  IBUFFX16_RVT U1 ( .A(\u_div/CryTmp[23][21] ), .Y(n1) );
  INVX2_RVT U2 ( .A(n1), .Y(n2) );
  INVX2_RVT U3 ( .A(n77), .Y(n78) );
  IBUFFX16_RVT U4 ( .A(\u_div/CryTmp[16][19] ), .Y(n77) );
  IBUFFX16_RVT U5 ( .A(\u_div/CryTmp[21][12] ), .Y(n3) );
  INVX4_RVT U6 ( .A(n3), .Y(n4) );
  IBUFFX2_RVT U7 ( .A(\u_div/CryTmp[18][14] ), .Y(n5) );
  IBUFFX4_RVT U8 ( .A(n5), .Y(n6) );
  IBUFFX16_RVT U9 ( .A(\u_div/CryTmp[18][20] ), .Y(n7) );
  INVX4_RVT U10 ( .A(n7), .Y(n8) );
  IBUFFX16_RVT U11 ( .A(\u_div/CryTmp[17][15] ), .Y(n9) );
  INVX4_RVT U12 ( .A(n9), .Y(n10) );
  IBUFFX16_RVT U13 ( .A(\u_div/CryTmp[24][12] ), .Y(n11) );
  INVX4_RVT U14 ( .A(n11), .Y(n12) );
  IBUFFX16_RVT U15 ( .A(\u_div/CryTmp[23][12] ), .Y(n13) );
  INVX4_RVT U16 ( .A(n13), .Y(n14) );
  IBUFFX16_RVT U17 ( .A(\u_div/CryTmp[24][17] ), .Y(n15) );
  INVX4_RVT U18 ( .A(n15), .Y(n16) );
  IBUFFX16_RVT U19 ( .A(\u_div/CryTmp[15][13] ), .Y(n17) );
  INVX4_RVT U20 ( .A(n17), .Y(n18) );
  IBUFFX16_RVT U21 ( .A(\u_div/CryTmp[18][12] ), .Y(n19) );
  INVX4_RVT U22 ( .A(n19), .Y(n20) );
  IBUFFX16_RVT U23 ( .A(\u_div/CryTmp[14][19] ), .Y(n21) );
  INVX4_RVT U24 ( .A(n21), .Y(n22) );
  IBUFFX16_RVT U25 ( .A(\u_div/CryTmp[18][13] ), .Y(n73) );
  INVX4_RVT U26 ( .A(n88), .Y(n23) );
  IBUFFX4_RVT U27 ( .A(n23), .Y(n24) );
  IBUFFX32_RVT U28 ( .A(n97), .Y(n25) );
  INVX0_RVT U29 ( .A(n25), .Y(n26) );
  INVX0_RVT U30 ( .A(n69), .Y(n27) );
  IBUFFX4_RVT U31 ( .A(n27), .Y(n28) );
  NOR2X2_RVT U32 ( .A1(\u_div/CryTmp[16][24] ), .A2(\u_div/PartRem[17][24] ), 
        .Y(n122) );
  INVX8_RVT U33 ( .A(n122), .Y(quotient[16]) );
  INVX4_RVT U34 ( .A(n117), .Y(n146) );
  INVX0_RVT U35 ( .A(n83), .Y(n84) );
  INVX1_RVT U36 ( .A(n344), .Y(\u_div/PartRem[18][21] ) );
  INVX1_RVT U37 ( .A(n52), .Y(n231) );
  INVX1_RVT U38 ( .A(\u_div/SumTmp[20][15] ), .Y(n475) );
  INVX1_RVT U39 ( .A(n116), .Y(n150) );
  INVX1_RVT U40 ( .A(n374), .Y(\u_div/PartRem[17][21] ) );
  INVX1_RVT U41 ( .A(n343), .Y(\u_div/PartRem[18][22] ) );
  INVX1_RVT U42 ( .A(n142), .Y(n141) );
  INVX1_RVT U43 ( .A(\u_div/CryTmp[24][24] ), .Y(\u_div/SumTmp[24][23] ) );
  INVX1_RVT U44 ( .A(\u_div/PartRem[21][23] ), .Y(n46) );
  INVX1_RVT U45 ( .A(\u_div/CryTmp[22][23] ), .Y(n81) );
  XOR2X1_RVT U46 ( .A1(\u_div/PartRem[18][23] ), .A2(\u_div/CryTmp[17][23] ), 
        .Y(\u_div/SumTmp[17][23] ) );
  OR2X1_RVT U47 ( .A1(n141), .A2(a[24]), .Y(\u_div/CryTmp[24][1] ) );
  MUX21X1_RVT U48 ( .A1(n208), .A2(n592), .S0(n146), .Y(n230) );
  INVX1_RVT U49 ( .A(n183), .Y(\u_div/PartRem[24][5] ) );
  MUX21X1_RVT U50 ( .A1(n207), .A2(n582), .S0(n146), .Y(n229) );
  INVX2_RVT U51 ( .A(n54), .Y(n55) );
  INVX1_RVT U52 ( .A(\u_div/SumTmp[20][2] ), .Y(n608) );
  MUX21X1_RVT U53 ( .A1(n206), .A2(n572), .S0(n146), .Y(n228) );
  MUX21X1_RVT U54 ( .A1(n205), .A2(n562), .S0(n146), .Y(n227) );
  INVX1_RVT U55 ( .A(\u_div/SumTmp[20][3] ), .Y(n600) );
  INVX1_RVT U56 ( .A(n48), .Y(n49) );
  INVX1_RVT U57 ( .A(\u_div/PartRem[17][1] ), .Y(n48) );
  INVX1_RVT U58 ( .A(n142), .Y(\u_div/CryTmp[23][1] ) );
  MUX21X1_RVT U59 ( .A1(n309), .A2(n621), .S0(quotient[18]), .Y(n334) );
  INVX1_RVT U60 ( .A(\u_div/SumTmp[18][2] ), .Y(n621) );
  MUX21X1_RVT U61 ( .A1(n204), .A2(n552), .S0(n146), .Y(n226) );
  INVX1_RVT U62 ( .A(n200), .Y(\u_div/PartRem[24][10] ) );
  MUX21X1_RVT U63 ( .A1(n202), .A2(n533), .S0(n146), .Y(n224) );
  MUX21X1_RVT U64 ( .A1(n201), .A2(n523), .S0(n146), .Y(n248) );
  INVX2_RVT U65 ( .A(n24), .Y(n89) );
  INVX1_RVT U66 ( .A(\u_div/SumTmp[20][9] ), .Y(n540) );
  INVX1_RVT U67 ( .A(n301), .Y(\u_div/PartRem[20][10] ) );
  MUX21X1_RVT U68 ( .A1(n221), .A2(n487), .S0(n146), .Y(n245) );
  INVX1_RVT U69 ( .A(n113), .Y(n105) );
  INVX1_RVT U70 ( .A(n113), .Y(n104) );
  INVX1_RVT U71 ( .A(n31), .Y(n45) );
  INVX1_RVT U72 ( .A(n30), .Y(n31) );
  INVX1_RVT U73 ( .A(n41), .Y(n148) );
  INVX1_RVT U74 ( .A(n113), .Y(n106) );
  INVX1_RVT U75 ( .A(n73), .Y(n74) );
  INVX1_RVT U76 ( .A(\u_div/SumTmp[18][12] ), .Y(n529) );
  INVX1_RVT U77 ( .A(n113), .Y(n107) );
  INVX1_RVT U78 ( .A(\u_div/SumTmp[20][16] ), .Y(n465) );
  IBUFFX4_RVT U79 ( .A(n126), .Y(n121) );
  INVX1_RVT U80 ( .A(n56), .Y(n57) );
  INVX1_RVT U81 ( .A(\u_div/CryTmp[18][17] ), .Y(n56) );
  INVX1_RVT U82 ( .A(n290), .Y(\u_div/PartRem[20][20] ) );
  MUX21X1_RVT U83 ( .A1(n266), .A2(n431), .S0(quotient[20]), .Y(n292) );
  INVX1_RVT U84 ( .A(\u_div/SumTmp[20][20] ), .Y(n368) );
  INVX1_RVT U85 ( .A(\u_div/SumTmp[21][22] ), .Y(n284) );
  INVX1_RVT U86 ( .A(\u_div/SumTmp[22][20] ), .Y(n311) );
  INVX1_RVT U87 ( .A(n101), .Y(n108) );
  INVX1_RVT U88 ( .A(n28), .Y(n70) );
  INVX1_RVT U89 ( .A(n315), .Y(\u_div/PartRem[19][21] ) );
  INVX1_RVT U90 ( .A(n345), .Y(\u_div/PartRem[18][20] ) );
  INVX1_RVT U91 ( .A(n408), .Y(\u_div/PartRem[16][19] ) );
  INVX1_RVT U92 ( .A(\u_div/SumTmp[20][21] ), .Y(n338) );
  INVX1_RVT U93 ( .A(\u_div/SumTmp[22][21] ), .Y(n285) );
  INVX2_RVT U94 ( .A(n90), .Y(n91) );
  INVX1_RVT U95 ( .A(n113), .Y(n114) );
  INVX2_RVT U96 ( .A(n36), .Y(n37) );
  INVX1_RVT U97 ( .A(n65), .Y(n66) );
  INVX1_RVT U98 ( .A(\u_div/CryTmp[16][23] ), .Y(n65) );
  INVX1_RVT U99 ( .A(n373), .Y(\u_div/PartRem[17][22] ) );
  NOR2X1_RVT U100 ( .A1(\u_div/PartRem[18][24] ), .A2(\u_div/CryTmp[17][24] ), 
        .Y(n123) );
  INVX1_RVT U101 ( .A(n99), .Y(n58) );
  OR2X1_RVT U102 ( .A1(\u_div/CryTmp[21][24] ), .A2(\u_div/PartRem[22][24] ), 
        .Y(quotient[21]) );
  INVX1_RVT U103 ( .A(\u_div/SumTmp[16][22] ), .Y(n427) );
  INVX1_RVT U104 ( .A(n53), .Y(n87) );
  DELLN2X2_RVT U105 ( .A(n26), .Y(n29) );
  INVX4_RVT U106 ( .A(n44), .Y(n30) );
  IBUFFX4_RVT U107 ( .A(\u_div/CryTmp[23][22] ), .Y(n32) );
  IBUFFX32_RVT U108 ( .A(n32), .Y(n33) );
  IBUFFX16_RVT U109 ( .A(\u_div/CryTmp[19][17] ), .Y(n34) );
  INVX4_RVT U110 ( .A(n34), .Y(n35) );
  IBUFFX4_RVT U111 ( .A(\u_div/CryTmp[19][23] ), .Y(n36) );
  INVX1_RVT U112 ( .A(n442), .Y(\u_div/PartRem[15][16] ) );
  INVX1_RVT U113 ( .A(n436), .Y(\u_div/PartRem[15][22] ) );
  OR2X2_RVT U114 ( .A1(\u_div/PartRem[16][24] ), .A2(\u_div/CryTmp[15][24] ), 
        .Y(quotient[15]) );
  INVX1_RVT U115 ( .A(\u_div/CryTmp[23][1] ), .Y(\u_div/SumTmp[18][0] ) );
  INVX1_RVT U116 ( .A(b[8]), .Y(\u_div/BInv[8] ) );
  INVX1_RVT U117 ( .A(b[7]), .Y(\u_div/BInv[7] ) );
  AND2X1_RVT U118 ( .A1(quotient[15]), .A2(\u_div/SumTmp[18][0] ), .Y(n39) );
  INVX1_RVT U119 ( .A(b[10]), .Y(\u_div/BInv[10] ) );
  AND2X1_RVT U120 ( .A1(n104), .A2(n127), .Y(n40) );
  INVX0_RVT U121 ( .A(n109), .Y(n113) );
  NOR2X1_RVT U122 ( .A1(n118), .A2(\u_div/PartRem[21][24] ), .Y(n41) );
  XNOR2X1_RVT U123 ( .A1(\u_div/CryTmp[19][10] ), .A2(n61), .Y(n43) );
  INVX1_RVT U124 ( .A(n292), .Y(\u_div/PartRem[20][19] ) );
  IBUFFX4_RVT U125 ( .A(\u_div/SumTmp[16][18] ), .Y(n481) );
  IBUFFX16_RVT U126 ( .A(\u_div/CryTmp[20][13] ), .Y(n44) );
  INVX2_RVT U127 ( .A(n46), .Y(n47) );
  INVX1_RVT U128 ( .A(n283), .Y(\u_div/PartRem[21][23] ) );
  IBUFFX4_RVT U129 ( .A(\u_div/PartRem[21][1] ), .Y(n50) );
  INVX4_RVT U130 ( .A(n50), .Y(n51) );
  MUX21X1_RVT U131 ( .A1(\u_div/SumTmp[22][1] ), .A2(n40), .S0(n117), .Y(n52)
         );
  MUX21X2_RVT U132 ( .A1(n222), .A2(n503), .S0(n146), .Y(n246) );
  MUX21X2_RVT U133 ( .A1(n223), .A2(n513), .S0(n146), .Y(n247) );
  MUX21X2_RVT U134 ( .A1(n203), .A2(n542), .S0(n146), .Y(n225) );
  IBUFFX4_RVT U135 ( .A(n293), .Y(\u_div/PartRem[20][18] ) );
  MUX21X2_RVT U136 ( .A1(n378), .A2(n481), .S0(quotient[16]), .Y(n408) );
  IBUFFX16_RVT U137 ( .A(quotient[15]), .Y(n53) );
  IBUFFX16_RVT U138 ( .A(\u_div/SumTmp[24][19] ), .Y(n287) );
  NOR2X2_RVT U139 ( .A1(\u_div/CryTmp[22][24] ), .A2(\u_div/PartRem[23][24] ), 
        .Y(n117) );
  IBUFFX16_RVT U140 ( .A(\u_div/SumTmp[23][22] ), .Y(n233) );
  INVX2_RVT U141 ( .A(a[24]), .Y(n594) );
  IBUFFX4_RVT U142 ( .A(n108), .Y(n109) );
  IBUFFX4_RVT U143 ( .A(\u_div/BInv[0] ), .Y(n142) );
  INVX1_RVT U144 ( .A(b[0]), .Y(\u_div/BInv[0] ) );
  INVX1_RVT U145 ( .A(\u_div/SumTmp[24][1] ), .Y(n584) );
  IBUFFX16_RVT U146 ( .A(\u_div/SumTmp[24][20] ), .Y(n260) );
  INVX0_RVT U147 ( .A(n291), .Y(\u_div/PartRem[20][1] ) );
  IBUFFX16_RVT U148 ( .A(\u_div/SumTmp[17][18] ), .Y(n472) );
  IBUFFX4_RVT U149 ( .A(\u_div/PartRem[20][2] ), .Y(n54) );
  INVX1_RVT U150 ( .A(n282), .Y(\u_div/PartRem[20][2] ) );
  IBUFFX4_RVT U151 ( .A(n98), .Y(n99) );
  IBUFFX4_RVT U152 ( .A(\u_div/PartRem[20][1] ), .Y(n59) );
  INVX4_RVT U153 ( .A(n59), .Y(n60) );
  IBUFFX4_RVT U154 ( .A(n108), .Y(n112) );
  XOR2X1_RVT U155 ( .A1(\u_div/PartRem[20][10] ), .A2(\u_div/BInv[10] ), .Y(
        n61) );
  NAND2X0_RVT U156 ( .A1(\u_div/PartRem[20][10] ), .A2(\u_div/CryTmp[19][10] ), 
        .Y(n62) );
  NAND2X0_RVT U157 ( .A1(\u_div/BInv[10] ), .A2(\u_div/CryTmp[19][10] ), .Y(
        n63) );
  NAND2X0_RVT U158 ( .A1(\u_div/BInv[10] ), .A2(\u_div/PartRem[20][10] ), .Y(
        n64) );
  NAND3X0_RVT U159 ( .A1(n62), .A2(n63), .A3(n64), .Y(\u_div/CryTmp[19][11] )
         );
  AND2X1_RVT U160 ( .A1(\u_div/CryTmp[23][23] ), .A2(\u_div/PartRem[24][23] ), 
        .Y(\u_div/CryTmp[23][24] ) );
  INVX16_RVT U161 ( .A(n238), .Y(n67) );
  IBUFFX16_RVT U162 ( .A(n67), .Y(n68) );
  IBUFFX16_RVT U163 ( .A(\u_div/CryTmp[24][22] ), .Y(n69) );
  IBUFFX16_RVT U164 ( .A(\u_div/CryTmp[16][17] ), .Y(n71) );
  INVX4_RVT U165 ( .A(n71), .Y(n72) );
  IBUFFX16_RVT U166 ( .A(\u_div/CryTmp[21][21] ), .Y(n75) );
  INVX4_RVT U167 ( .A(n75), .Y(n76) );
  IBUFFX16_RVT U168 ( .A(\u_div/CryTmp[24][21] ), .Y(n79) );
  INVX4_RVT U169 ( .A(n79), .Y(n80) );
  IBUFFX4_RVT U170 ( .A(n81), .Y(n82) );
  IBUFFX16_RVT U171 ( .A(\u_div/CryTmp[15][18] ), .Y(n83) );
  IBUFFX16_RVT U172 ( .A(\u_div/CryTmp[17][21] ), .Y(n85) );
  INVX4_RVT U173 ( .A(n85), .Y(n86) );
  IBUFFX16_RVT U174 ( .A(\u_div/CryTmp[22][13] ), .Y(n88) );
  IBUFFX16_RVT U175 ( .A(\u_div/CryTmp[22][22] ), .Y(n90) );
  IBUFFX16_RVT U176 ( .A(\u_div/CryTmp[14][22] ), .Y(n92) );
  INVX4_RVT U177 ( .A(n92), .Y(n93) );
  IBUFFX16_RVT U178 ( .A(\u_div/CryTmp[20][22] ), .Y(n94) );
  INVX4_RVT U179 ( .A(n94), .Y(n95) );
  NOR2X2_RVT U180 ( .A1(\u_div/CryTmp[18][24] ), .A2(\u_div/PartRem[19][24] ), 
        .Y(n119) );
  INVX2_RVT U181 ( .A(n336), .Y(\u_div/PartRem[19][23] ) );
  INVX32_RVT U182 ( .A(\u_div/CryTmp[18][23] ), .Y(n96) );
  IBUFFX16_RVT U183 ( .A(n96), .Y(n97) );
  IBUFFX4_RVT U184 ( .A(n150), .Y(n98) );
  INVX2_RVT U185 ( .A(n98), .Y(n100) );
  INVX0_RVT U186 ( .A(n145), .Y(n101) );
  NBUFFX2_RVT U187 ( .A(n145), .Y(n102) );
  INVX1_RVT U188 ( .A(n102), .Y(n103) );
  INVX1_RVT U189 ( .A(n108), .Y(n110) );
  INVX1_RVT U190 ( .A(n108), .Y(n111) );
  INVX1_RVT U191 ( .A(n113), .Y(quotient[23]) );
  OR2X1_RVT U192 ( .A1(\u_div/CryTmp[23][24] ), .A2(\u_div/PartRem[24][24] ), 
        .Y(n629) );
  IBUFFX4_RVT U193 ( .A(n629), .Y(n145) );
  INVX1_RVT U194 ( .A(n307), .Y(\u_div/PartRem[19][4] ) );
  INVX1_RVT U195 ( .A(n264), .Y(\u_div/PartRem[21][1] ) );
  INVX1_RVT U196 ( .A(n308), .Y(\u_div/PartRem[19][3] ) );
  INVX0_RVT U197 ( .A(b[12]), .Y(\u_div/BInv[12] ) );
  INVX0_RVT U198 ( .A(b[11]), .Y(\u_div/BInv[11] ) );
  INVX0_RVT U199 ( .A(b[21]), .Y(\u_div/BInv[21] ) );
  INVX0_RVT U200 ( .A(b[20]), .Y(\u_div/BInv[20] ) );
  INVX0_RVT U201 ( .A(b[19]), .Y(\u_div/BInv[19] ) );
  INVX0_RVT U202 ( .A(b[18]), .Y(\u_div/BInv[18] ) );
  INVX0_RVT U203 ( .A(b[16]), .Y(\u_div/BInv[16] ) );
  INVX0_RVT U204 ( .A(b[17]), .Y(\u_div/BInv[17] ) );
  INVX4_RVT U205 ( .A(n123), .Y(n154) );
  INVX4_RVT U206 ( .A(n119), .Y(n152) );
  INVX0_RVT U207 ( .A(n119), .Y(quotient[18]) );
  INVX0_RVT U208 ( .A(n123), .Y(quotient[17]) );
  INVX0_RVT U209 ( .A(n58), .Y(quotient[19]) );
  INVX1_RVT U210 ( .A(n281), .Y(\u_div/PartRem[20][3] ) );
  INVX0_RVT U211 ( .A(\u_div/CryTmp[23][1] ), .Y(\u_div/SumTmp[20][0] ) );
  INVX0_RVT U212 ( .A(n623), .Y(n130) );
  INVX0_RVT U213 ( .A(\u_div/CryTmp[23][1] ), .Y(\u_div/SumTmp[19][0] ) );
  INVX0_RVT U214 ( .A(n628), .Y(n131) );
  INVX0_RVT U215 ( .A(\u_div/CryTmp[23][1] ), .Y(\u_div/SumTmp[21][0] ) );
  INVX0_RVT U216 ( .A(n617), .Y(n129) );
  AND2X1_RVT U217 ( .A1(n82), .A2(\u_div/PartRem[23][23] ), .Y(
        \u_div/CryTmp[22][24] ) );
  AND2X1_RVT U218 ( .A1(n37), .A2(n124), .Y(\u_div/CryTmp[19][24] ) );
  AND2X1_RVT U219 ( .A1(\u_div/CryTmp[21][23] ), .A2(\u_div/PartRem[22][23] ), 
        .Y(\u_div/CryTmp[21][24] ) );
  INVX1_RVT U220 ( .A(n365), .Y(\u_div/PartRem[18][23] ) );
  INVX1_RVT U221 ( .A(\u_div/SumTmp[18][22] ), .Y(n366) );
  INVX1_RVT U222 ( .A(n256), .Y(\u_div/PartRem[21][2] ) );
  INVX0_RVT U223 ( .A(\u_div/CryTmp[23][1] ), .Y(\u_div/SumTmp[22][0] ) );
  INVX0_RVT U224 ( .A(n610), .Y(n128) );
  INVX0_RVT U225 ( .A(n144), .Y(n120) );
  INVX1_RVT U226 ( .A(n328), .Y(\u_div/PartRem[18][9] ) );
  INVX1_RVT U227 ( .A(n276), .Y(\u_div/PartRem[20][8] ) );
  INVX1_RVT U228 ( .A(n303), .Y(\u_div/PartRem[19][8] ) );
  INVX1_RVT U229 ( .A(n277), .Y(\u_div/PartRem[20][7] ) );
  INVX1_RVT U230 ( .A(n394), .Y(\u_div/PartRem[16][2] ) );
  INVX1_RVT U231 ( .A(n393), .Y(\u_div/PartRem[16][3] ) );
  INVX0_RVT U232 ( .A(\u_div/CryTmp[23][1] ), .Y(\u_div/SumTmp[23][0] ) );
  INVX0_RVT U233 ( .A(n602), .Y(n127) );
  INVX1_RVT U234 ( .A(n392), .Y(\u_div/PartRem[16][4] ) );
  INVX1_RVT U235 ( .A(n445), .Y(\u_div/PartRem[15][13] ) );
  INVX1_RVT U236 ( .A(\u_div/SumTmp[15][12] ), .Y(n555) );
  INVX1_RVT U237 ( .A(n443), .Y(\u_div/PartRem[15][15] ) );
  INVX1_RVT U238 ( .A(\u_div/SumTmp[15][14] ), .Y(n536) );
  INVX1_RVT U239 ( .A(n232), .Y(\u_div/PartRem[23][23] ) );
  AND2X1_RVT U240 ( .A1(\u_div/CryTmp[17][23] ), .A2(\u_div/PartRem[18][23] ), 
        .Y(\u_div/CryTmp[17][24] ) );
  NOR2X0_RVT U241 ( .A1(\u_div/CryTmp[19][24] ), .A2(\u_div/PartRem[20][24] ), 
        .Y(n116) );
  AND2X1_RVT U242 ( .A1(n66), .A2(\u_div/PartRem[17][23] ), .Y(
        \u_div/CryTmp[16][24] ) );
  AND2X1_RVT U243 ( .A1(\u_div/CryTmp[15][23] ), .A2(\u_div/PartRem[16][23] ), 
        .Y(\u_div/CryTmp[15][24] ) );
  AND2X1_RVT U244 ( .A1(\u_div/CryTmp[20][23] ), .A2(n47), .Y(n118) );
  MUX21X1_RVT U245 ( .A1(\u_div/PartRem[21][22] ), .A2(\u_div/SumTmp[20][22] ), 
        .S0(quotient[20]), .Y(n124) );
  INVX1_RVT U246 ( .A(n426), .Y(\u_div/PartRem[16][23] ) );
  INVX1_RVT U247 ( .A(n257), .Y(\u_div/PartRem[22][23] ) );
  INVX1_RVT U248 ( .A(\u_div/SumTmp[22][22] ), .Y(n258) );
  INVX1_RVT U249 ( .A(\u_div/SumTmp[19][22] ), .Y(n337) );
  INVX1_RVT U250 ( .A(n395), .Y(\u_div/PartRem[17][23] ) );
  INVX1_RVT U251 ( .A(\u_div/SumTmp[17][22] ), .Y(n396) );
  INVX1_RVT U252 ( .A(n187), .Y(\u_div/PartRem[24][22] ) );
  INVX1_RVT U253 ( .A(n211), .Y(\u_div/PartRem[23][22] ) );
  INVX1_RVT U254 ( .A(n235), .Y(\u_div/PartRem[22][22] ) );
  INVX1_RVT U255 ( .A(n404), .Y(\u_div/PartRem[16][22] ) );
  INVX1_RVT U256 ( .A(n298), .Y(\u_div/PartRem[20][13] ) );
  INVX1_RVT U257 ( .A(n297), .Y(\u_div/PartRem[20][14] ) );
  INVX1_RVT U258 ( .A(n296), .Y(\u_div/PartRem[20][15] ) );
  INVX1_RVT U259 ( .A(n383), .Y(\u_div/PartRem[17][13] ) );
  INVX1_RVT U260 ( .A(n414), .Y(\u_div/PartRem[16][13] ) );
  INVX1_RVT U261 ( .A(n413), .Y(\u_div/PartRem[16][14] ) );
  INVX1_RVT U262 ( .A(n412), .Y(\u_div/PartRem[16][15] ) );
  INVX1_RVT U263 ( .A(n444), .Y(\u_div/PartRem[15][14] ) );
  INVX1_RVT U264 ( .A(n326), .Y(\u_div/PartRem[19][11] ) );
  INVX1_RVT U265 ( .A(n188), .Y(\u_div/PartRem[24][21] ) );
  INVX1_RVT U266 ( .A(n189), .Y(\u_div/PartRem[24][20] ) );
  INVX1_RVT U267 ( .A(n191), .Y(\u_div/PartRem[24][19] ) );
  INVX1_RVT U268 ( .A(n192), .Y(\u_div/PartRem[24][18] ) );
  INVX1_RVT U269 ( .A(n193), .Y(\u_div/PartRem[24][17] ) );
  INVX1_RVT U270 ( .A(n266), .Y(\u_div/PartRem[21][18] ) );
  INVX1_RVT U271 ( .A(n265), .Y(\u_div/PartRem[21][19] ) );
  INVX1_RVT U272 ( .A(n262), .Y(\u_div/PartRem[21][21] ) );
  INVX1_RVT U273 ( .A(n295), .Y(\u_div/PartRem[20][16] ) );
  INVX1_RVT U274 ( .A(n320), .Y(\u_div/PartRem[19][17] ) );
  INVX1_RVT U275 ( .A(n319), .Y(\u_div/PartRem[19][18] ) );
  INVX1_RVT U276 ( .A(n354), .Y(\u_div/PartRem[18][12] ) );
  INVX1_RVT U277 ( .A(n384), .Y(\u_div/PartRem[17][12] ) );
  INVX1_RVT U278 ( .A(n415), .Y(\u_div/PartRem[16][12] ) );
  INVX1_RVT U279 ( .A(n411), .Y(\u_div/PartRem[16][16] ) );
  INVX1_RVT U280 ( .A(n410), .Y(\u_div/PartRem[16][17] ) );
  INVX1_RVT U281 ( .A(n409), .Y(\u_div/PartRem[16][18] ) );
  INVX1_RVT U282 ( .A(n406), .Y(\u_div/PartRem[16][20] ) );
  INVX1_RVT U283 ( .A(n405), .Y(\u_div/PartRem[16][21] ) );
  INVX1_RVT U284 ( .A(n446), .Y(\u_div/PartRem[15][12] ) );
  INVX1_RVT U285 ( .A(n356), .Y(\u_div/PartRem[18][10] ) );
  INVX1_RVT U286 ( .A(n386), .Y(\u_div/PartRem[17][10] ) );
  INVX1_RVT U287 ( .A(n355), .Y(\u_div/PartRem[18][11] ) );
  INVX1_RVT U288 ( .A(n385), .Y(\u_div/PartRem[17][11] ) );
  INVX1_RVT U289 ( .A(n416), .Y(\u_div/PartRem[16][11] ) );
  INVX1_RVT U290 ( .A(n327), .Y(\u_div/PartRem[19][10] ) );
  INVX1_RVT U291 ( .A(n209), .Y(\u_div/PartRem[24][23] ) );
  INVX1_RVT U292 ( .A(\u_div/SumTmp[24][22] ), .Y(n210) );
  INVX1_RVT U293 ( .A(n424), .Y(\u_div/PartRem[15][3] ) );
  INVX1_RVT U294 ( .A(n422), .Y(\u_div/PartRem[15][5] ) );
  INVX1_RVT U295 ( .A(n41), .Y(quotient[20]) );
  INVX1_RVT U296 ( .A(n117), .Y(quotient[22]) );
  INVX1_RVT U297 ( .A(\u_div/SumTmp[24][23] ), .Y(n144) );
  INVX1_RVT U298 ( .A(n121), .Y(n143) );
  INVX1_RVT U299 ( .A(\u_div/SumTmp[24][23] ), .Y(n126) );
  OR2X1_RVT U300 ( .A1(n120), .A2(n121), .Y(\u_div/PartRem[24][24] ) );
  INVX1_RVT U301 ( .A(n255), .Y(\u_div/PartRem[21][3] ) );
  INVX1_RVT U302 ( .A(n280), .Y(\u_div/PartRem[20][4] ) );
  INVX1_RVT U303 ( .A(n407), .Y(\u_div/PartRem[16][1] ) );
  INVX1_RVT U304 ( .A(n306), .Y(\u_div/PartRem[19][5] ) );
  INVX1_RVT U305 ( .A(n201), .Y(\u_div/PartRem[23][9] ) );
  INVX1_RVT U306 ( .A(n202), .Y(\u_div/PartRem[23][8] ) );
  INVX1_RVT U307 ( .A(n203), .Y(\u_div/PartRem[23][7] ) );
  INVX1_RVT U308 ( .A(n204), .Y(\u_div/PartRem[23][6] ) );
  INVX1_RVT U309 ( .A(n205), .Y(\u_div/PartRem[23][5] ) );
  INVX1_RVT U310 ( .A(n206), .Y(\u_div/PartRem[23][4] ) );
  INVX1_RVT U311 ( .A(n207), .Y(\u_div/PartRem[23][3] ) );
  INVX1_RVT U312 ( .A(n208), .Y(\u_div/PartRem[23][2] ) );
  INVX0_RVT U313 ( .A(n224), .Y(\u_div/PartRem[22][9] ) );
  INVX1_RVT U314 ( .A(n225), .Y(\u_div/PartRem[22][8] ) );
  INVX1_RVT U315 ( .A(n226), .Y(\u_div/PartRem[22][7] ) );
  INVX1_RVT U316 ( .A(n227), .Y(\u_div/PartRem[22][6] ) );
  INVX1_RVT U317 ( .A(n228), .Y(\u_div/PartRem[22][5] ) );
  INVX1_RVT U318 ( .A(n229), .Y(\u_div/PartRem[22][4] ) );
  INVX1_RVT U319 ( .A(n230), .Y(\u_div/PartRem[22][3] ) );
  INVX1_RVT U320 ( .A(n254), .Y(\u_div/PartRem[21][4] ) );
  INVX1_RVT U321 ( .A(n249), .Y(\u_div/PartRem[21][9] ) );
  INVX1_RVT U322 ( .A(n250), .Y(\u_div/PartRem[21][8] ) );
  INVX1_RVT U323 ( .A(n251), .Y(\u_div/PartRem[21][7] ) );
  INVX1_RVT U324 ( .A(n252), .Y(\u_div/PartRem[21][6] ) );
  INVX1_RVT U325 ( .A(n253), .Y(\u_div/PartRem[21][5] ) );
  INVX1_RVT U326 ( .A(n363), .Y(\u_div/PartRem[17][3] ) );
  INVX1_RVT U327 ( .A(n364), .Y(\u_div/PartRem[17][2] ) );
  INVX1_RVT U328 ( .A(n279), .Y(\u_div/PartRem[20][5] ) );
  INVX1_RVT U329 ( .A(n335), .Y(\u_div/PartRem[18][2] ) );
  INVX1_RVT U330 ( .A(n357), .Y(\u_div/PartRem[17][9] ) );
  INVX1_RVT U331 ( .A(n346), .Y(\u_div/PartRem[18][1] ) );
  INVX1_RVT U332 ( .A(n388), .Y(\u_div/PartRem[16][8] ) );
  INVX1_RVT U333 ( .A(n305), .Y(\u_div/PartRem[19][6] ) );
  INVX1_RVT U334 ( .A(n425), .Y(\u_div/PartRem[15][2] ) );
  INVX1_RVT U335 ( .A(n423), .Y(\u_div/PartRem[15][4] ) );
  INVX1_RVT U336 ( .A(n304), .Y(\u_div/PartRem[19][7] ) );
  INVX1_RVT U337 ( .A(n302), .Y(\u_div/PartRem[19][9] ) );
  INVX1_RVT U338 ( .A(n278), .Y(\u_div/PartRem[20][6] ) );
  INVX1_RVT U339 ( .A(n275), .Y(\u_div/PartRem[20][9] ) );
  INVX1_RVT U340 ( .A(n376), .Y(\u_div/PartRem[17][1] ) );
  INVX1_RVT U341 ( .A(n387), .Y(\u_div/PartRem[16][9] ) );
  AND2X1_RVT U342 ( .A1(n29), .A2(\u_div/PartRem[19][23] ), .Y(
        \u_div/CryTmp[18][24] ) );
  INVX1_RVT U343 ( .A(n419), .Y(\u_div/PartRem[15][8] ) );
  INVX1_RVT U344 ( .A(n441), .Y(\u_div/PartRem[15][17] ) );
  INVX1_RVT U345 ( .A(n439), .Y(\u_div/PartRem[15][19] ) );
  INVX1_RVT U346 ( .A(n437), .Y(\u_div/PartRem[15][21] ) );
  XOR2X1_RVT U347 ( .A1(\u_div/PartRem[17][23] ), .A2(n66), .Y(
        \u_div/SumTmp[16][23] ) );
  XOR2X1_RVT U348 ( .A1(\u_div/PartRem[16][23] ), .A2(\u_div/CryTmp[15][23] ), 
        .Y(\u_div/SumTmp[15][23] ) );
  XOR2X1_RVT U349 ( .A1(\u_div/PartRem[19][23] ), .A2(n29), .Y(
        \u_div/SumTmp[18][23] ) );
  INVX1_RVT U350 ( .A(n449), .Y(\u_div/PartRem[15][23] ) );
  INVX1_RVT U351 ( .A(n317), .Y(\u_div/PartRem[19][1] ) );
  INVX1_RVT U352 ( .A(n309), .Y(\u_div/PartRem[19][2] ) );
  XOR2X1_RVT U353 ( .A1(n124), .A2(n37), .Y(\u_div/SumTmp[19][23] ) );
  XOR2X1_RVT U354 ( .A1(n47), .A2(\u_div/CryTmp[20][23] ), .Y(
        \u_div/SumTmp[20][23] ) );
  XOR2X1_RVT U355 ( .A1(\u_div/PartRem[22][23] ), .A2(\u_div/CryTmp[21][23] ), 
        .Y(\u_div/SumTmp[21][23] ) );
  INVX1_RVT U356 ( .A(n68), .Y(\u_div/PartRem[22][1] ) );
  MUX21X1_RVT U357 ( .A1(n236), .A2(n310), .S0(quotient[21]), .Y(n261) );
  XOR2X1_RVT U358 ( .A1(\u_div/PartRem[23][23] ), .A2(n82), .Y(
        \u_div/SumTmp[22][23] ) );
  INVX1_RVT U359 ( .A(n186), .Y(\u_div/PartRem[24][2] ) );
  INVX1_RVT U360 ( .A(n185), .Y(\u_div/PartRem[24][3] ) );
  INVX1_RVT U361 ( .A(n184), .Y(\u_div/PartRem[24][4] ) );
  INVX1_RVT U362 ( .A(n182), .Y(\u_div/PartRem[24][6] ) );
  INVX1_RVT U363 ( .A(n181), .Y(\u_div/PartRem[24][7] ) );
  INVX1_RVT U364 ( .A(n180), .Y(\u_div/PartRem[24][8] ) );
  INVX1_RVT U365 ( .A(n179), .Y(\u_div/PartRem[24][9] ) );
  XOR2X1_RVT U366 ( .A1(\u_div/PartRem[24][23] ), .A2(\u_div/CryTmp[23][23] ), 
        .Y(\u_div/SumTmp[23][23] ) );
  INVX1_RVT U367 ( .A(n212), .Y(\u_div/PartRem[23][21] ) );
  INVX1_RVT U368 ( .A(n213), .Y(\u_div/PartRem[23][20] ) );
  INVX1_RVT U369 ( .A(n214), .Y(\u_div/PartRem[23][19] ) );
  INVX1_RVT U370 ( .A(n215), .Y(\u_div/PartRem[23][18] ) );
  INVX1_RVT U371 ( .A(n239), .Y(\u_div/PartRem[22][19] ) );
  INVX1_RVT U372 ( .A(n236), .Y(\u_div/PartRem[22][21] ) );
  INVX1_RVT U373 ( .A(n263), .Y(\u_div/PartRem[21][20] ) );
  INVX1_RVT U374 ( .A(n289), .Y(\u_div/PartRem[20][21] ) );
  INVX1_RVT U375 ( .A(n314), .Y(\u_div/PartRem[19][22] ) );
  INVX1_RVT U376 ( .A(n219), .Y(\u_div/PartRem[23][14] ) );
  INVX1_RVT U377 ( .A(n220), .Y(\u_div/PartRem[23][13] ) );
  INVX1_RVT U378 ( .A(n221), .Y(\u_div/PartRem[23][12] ) );
  INVX1_RVT U379 ( .A(n222), .Y(\u_div/PartRem[23][11] ) );
  INVX1_RVT U380 ( .A(n223), .Y(\u_div/PartRem[23][10] ) );
  INVX0_RVT U381 ( .A(n244), .Y(\u_div/PartRem[22][14] ) );
  INVX1_RVT U382 ( .A(n245), .Y(\u_div/PartRem[22][13] ) );
  INVX1_RVT U383 ( .A(n246), .Y(\u_div/PartRem[22][12] ) );
  INVX1_RVT U384 ( .A(n247), .Y(\u_div/PartRem[22][11] ) );
  INVX1_RVT U385 ( .A(n248), .Y(\u_div/PartRem[22][10] ) );
  INVX1_RVT U386 ( .A(n269), .Y(\u_div/PartRem[21][15] ) );
  INVX1_RVT U387 ( .A(n270), .Y(\u_div/PartRem[21][14] ) );
  INVX1_RVT U388 ( .A(n271), .Y(\u_div/PartRem[21][13] ) );
  INVX1_RVT U389 ( .A(n272), .Y(\u_div/PartRem[21][12] ) );
  INVX1_RVT U390 ( .A(n273), .Y(\u_div/PartRem[21][11] ) );
  INVX1_RVT U391 ( .A(n274), .Y(\u_div/PartRem[21][10] ) );
  INVX1_RVT U392 ( .A(n242), .Y(\u_div/PartRem[22][16] ) );
  INVX1_RVT U393 ( .A(n380), .Y(\u_div/PartRem[17][16] ) );
  INVX1_RVT U394 ( .A(n381), .Y(\u_div/PartRem[17][15] ) );
  INVX1_RVT U395 ( .A(n382), .Y(\u_div/PartRem[17][14] ) );
  INVX1_RVT U396 ( .A(n375), .Y(\u_div/PartRem[17][20] ) );
  INVX1_RVT U397 ( .A(n377), .Y(\u_div/PartRem[17][19] ) );
  INVX1_RVT U398 ( .A(n378), .Y(\u_div/PartRem[17][18] ) );
  INVX1_RVT U399 ( .A(n379), .Y(\u_div/PartRem[17][17] ) );
  INVX1_RVT U400 ( .A(n351), .Y(\u_div/PartRem[18][15] ) );
  INVX1_RVT U401 ( .A(n353), .Y(\u_div/PartRem[18][13] ) );
  INVX1_RVT U402 ( .A(n352), .Y(\u_div/PartRem[18][14] ) );
  INVX1_RVT U403 ( .A(n347), .Y(\u_div/PartRem[18][19] ) );
  INVX1_RVT U404 ( .A(n348), .Y(\u_div/PartRem[18][18] ) );
  INVX1_RVT U405 ( .A(n349), .Y(\u_div/PartRem[18][17] ) );
  INVX1_RVT U406 ( .A(n350), .Y(\u_div/PartRem[18][16] ) );
  INVX1_RVT U407 ( .A(n318), .Y(\u_div/PartRem[19][19] ) );
  INVX1_RVT U408 ( .A(n440), .Y(\u_div/PartRem[15][18] ) );
  INVX1_RVT U409 ( .A(n325), .Y(\u_div/PartRem[19][12] ) );
  INVX1_RVT U410 ( .A(n324), .Y(\u_div/PartRem[19][13] ) );
  INVX1_RVT U411 ( .A(n323), .Y(\u_div/PartRem[19][14] ) );
  INVX1_RVT U412 ( .A(n300), .Y(\u_div/PartRem[20][11] ) );
  INVX1_RVT U413 ( .A(n299), .Y(\u_div/PartRem[20][12] ) );
  INVX1_RVT U414 ( .A(n438), .Y(\u_div/PartRem[15][20] ) );
  INVX1_RVT U415 ( .A(n294), .Y(\u_div/PartRem[20][17] ) );
  INVX1_RVT U416 ( .A(b[9]), .Y(n132) );
  INVX1_RVT U417 ( .A(b[6]), .Y(n133) );
  INVX1_RVT U418 ( .A(b[5]), .Y(n134) );
  INVX1_RVT U419 ( .A(b[4]), .Y(n135) );
  INVX1_RVT U420 ( .A(b[3]), .Y(n136) );
  INVX1_RVT U421 ( .A(b[2]), .Y(n137) );
  INVX1_RVT U422 ( .A(b[1]), .Y(n139) );
  INVX1_RVT U423 ( .A(n190), .Y(\u_div/PartRem[24][1] ) );
  INVX1_RVT U424 ( .A(n197), .Y(\u_div/PartRem[24][13] ) );
  INVX1_RVT U425 ( .A(n199), .Y(\u_div/PartRem[24][11] ) );
  INVX1_RVT U426 ( .A(n198), .Y(\u_div/PartRem[24][12] ) );
  INVX1_RVT U427 ( .A(n196), .Y(\u_div/PartRem[24][14] ) );
  INVX1_RVT U428 ( .A(b[1]), .Y(n140) );
  INVX1_RVT U429 ( .A(b[2]), .Y(n138) );
  INVX1_RVT U430 ( .A(b[15]), .Y(\u_div/BInv[15] ) );
  INVX1_RVT U431 ( .A(b[14]), .Y(\u_div/BInv[14] ) );
  INVX1_RVT U432 ( .A(b[13]), .Y(\u_div/BInv[13] ) );
  OR2X1_RVT U433 ( .A1(\u_div/CryTmp[14][24] ), .A2(\u_div/PartRem[15][24] ), 
        .Y(quotient[14]) );
  AND2X1_RVT U434 ( .A1(\u_div/PartRem[15][23] ), .A2(\u_div/CryTmp[14][23] ), 
        .Y(\u_div/CryTmp[14][24] ) );
  INVX1_RVT U435 ( .A(b[6]), .Y(\u_div/BInv[6] ) );
  INVX1_RVT U436 ( .A(b[5]), .Y(\u_div/BInv[5] ) );
  INVX1_RVT U437 ( .A(b[4]), .Y(\u_div/BInv[4] ) );
  INVX1_RVT U438 ( .A(b[3]), .Y(\u_div/BInv[3] ) );
  XNOR2X1_RVT U439 ( .A1(n594), .A2(n141), .Y(n125) );
  NAND2X0_RVT U440 ( .A1(n146), .A2(n128), .Y(n238) );
  NAND2X0_RVT U441 ( .A1(quotient[21]), .A2(n129), .Y(n264) );
  NAND2X0_RVT U442 ( .A1(n148), .A2(n130), .Y(n291) );
  NAND2X0_RVT U443 ( .A1(n99), .A2(n131), .Y(n317) );
  NAND2X0_RVT U444 ( .A1(n152), .A2(\u_div/SumTmp[18][0] ), .Y(n346) );
  NAND2X0_RVT U445 ( .A1(n154), .A2(\u_div/SumTmp[18][0] ), .Y(n376) );
  NAND2X0_RVT U446 ( .A1(quotient[16]), .A2(\u_div/SumTmp[18][0] ), .Y(n407)
         );
  INVX1_RVT U447 ( .A(n329), .Y(\u_div/PartRem[18][8] ) );
  INVX1_RVT U448 ( .A(n288), .Y(\u_div/PartRem[20][22] ) );
  INVX1_RVT U449 ( .A(b[22]), .Y(\u_div/BInv[22] ) );
  INVX1_RVT U450 ( .A(n447), .Y(\u_div/PartRem[15][11] ) );
  INVX1_RVT U451 ( .A(n417), .Y(\u_div/PartRem[16][10] ) );
  INVX1_RVT U452 ( .A(n358), .Y(\u_div/PartRem[17][8] ) );
  INVX1_RVT U453 ( .A(n330), .Y(\u_div/PartRem[18][7] ) );
  INVX1_RVT U454 ( .A(n321), .Y(\u_div/PartRem[19][16] ) );
  INVX1_RVT U455 ( .A(n261), .Y(\u_div/PartRem[21][22] ) );
  INVX1_RVT U456 ( .A(n237), .Y(\u_div/PartRem[22][20] ) );
  INVX1_RVT U457 ( .A(n216), .Y(\u_div/PartRem[23][17] ) );
  INVX1_RVT U458 ( .A(n448), .Y(\u_div/PartRem[15][10] ) );
  INVX1_RVT U459 ( .A(n331), .Y(\u_div/PartRem[18][6] ) );
  INVX1_RVT U460 ( .A(n240), .Y(\u_div/PartRem[22][18] ) );
  INVX1_RVT U461 ( .A(n217), .Y(\u_div/PartRem[23][16] ) );
  INVX1_RVT U462 ( .A(n389), .Y(\u_div/PartRem[16][7] ) );
  INVX1_RVT U463 ( .A(n359), .Y(\u_div/PartRem[17][7] ) );
  INVX1_RVT U464 ( .A(n332), .Y(\u_div/PartRem[18][5] ) );
  INVX1_RVT U465 ( .A(n322), .Y(\u_div/PartRem[19][15] ) );
  INVX1_RVT U466 ( .A(n243), .Y(\u_div/PartRem[22][15] ) );
  INVX1_RVT U467 ( .A(n390), .Y(\u_div/PartRem[16][6] ) );
  INVX1_RVT U468 ( .A(n241), .Y(\u_div/PartRem[22][17] ) );
  INVX1_RVT U469 ( .A(n418), .Y(\u_div/PartRem[15][9] ) );
  INVX1_RVT U470 ( .A(n360), .Y(\u_div/PartRem[17][6] ) );
  INVX1_RVT U471 ( .A(n333), .Y(\u_div/PartRem[18][4] ) );
  INVX1_RVT U472 ( .A(n316), .Y(\u_div/PartRem[19][20] ) );
  INVX1_RVT U473 ( .A(n194), .Y(\u_div/PartRem[24][16] ) );
  INVX1_RVT U474 ( .A(n195), .Y(\u_div/PartRem[24][15] ) );
  INVX1_RVT U475 ( .A(n420), .Y(\u_div/PartRem[15][7] ) );
  INVX1_RVT U476 ( .A(n391), .Y(\u_div/PartRem[16][5] ) );
  INVX1_RVT U477 ( .A(n362), .Y(\u_div/PartRem[17][4] ) );
  INVX1_RVT U478 ( .A(n361), .Y(\u_div/PartRem[17][5] ) );
  INVX1_RVT U479 ( .A(n334), .Y(\u_div/PartRem[18][3] ) );
  INVX1_RVT U480 ( .A(n267), .Y(\u_div/PartRem[21][17] ) );
  INVX1_RVT U481 ( .A(n218), .Y(\u_div/PartRem[23][15] ) );
  INVX1_RVT U482 ( .A(n421), .Y(\u_div/PartRem[15][6] ) );
  MUX21X1_RVT U483 ( .A1(\u_div/PartRem[24][23] ), .A2(\u_div/SumTmp[23][23] ), 
        .S0(n114), .Y(\u_div/PartRem[23][24] ) );
  MUX21X1_RVT U484 ( .A1(n165), .A2(n210), .S0(n144), .Y(n209) );
  INVX0_RVT U485 ( .A(a[46]), .Y(n165) );
  MUX21X1_RVT U486 ( .A1(\u_div/PartRem[23][23] ), .A2(\u_div/SumTmp[22][23] ), 
        .S0(quotient[22]), .Y(\u_div/PartRem[22][24] ) );
  MUX21X1_RVT U487 ( .A1(n187), .A2(n233), .S0(n112), .Y(n232) );
  MUX21X1_RVT U488 ( .A1(n166), .A2(n234), .S0(n144), .Y(n187) );
  INVX0_RVT U489 ( .A(\u_div/SumTmp[24][21] ), .Y(n234) );
  INVX0_RVT U490 ( .A(a[45]), .Y(n166) );
  MUX21X1_RVT U491 ( .A1(\u_div/PartRem[22][23] ), .A2(\u_div/SumTmp[21][23] ), 
        .S0(quotient[21]), .Y(\u_div/PartRem[21][24] ) );
  MUX21X1_RVT U492 ( .A1(n211), .A2(n258), .S0(quotient[22]), .Y(n257) );
  MUX21X1_RVT U493 ( .A1(n188), .A2(n259), .S0(n111), .Y(n211) );
  INVX0_RVT U494 ( .A(\u_div/SumTmp[23][21] ), .Y(n259) );
  MUX21X1_RVT U495 ( .A1(n167), .A2(n260), .S0(n144), .Y(n188) );
  INVX0_RVT U496 ( .A(a[44]), .Y(n167) );
  IBUFFX16_RVT U497 ( .A(n268), .Y(\u_div/PartRem[21][16] ) );
  MUX21X1_RVT U498 ( .A1(n47), .A2(\u_div/SumTmp[20][23] ), .S0(quotient[20]), 
        .Y(\u_div/PartRem[20][24] ) );
  MUX21X1_RVT U499 ( .A1(n235), .A2(n284), .S0(quotient[21]), .Y(n283) );
  MUX21X1_RVT U500 ( .A1(n212), .A2(n285), .S0(quotient[22]), .Y(n235) );
  MUX21X1_RVT U501 ( .A1(n189), .A2(n286), .S0(n110), .Y(n212) );
  INVX0_RVT U502 ( .A(\u_div/SumTmp[23][20] ), .Y(n286) );
  MUX21X1_RVT U503 ( .A1(n169), .A2(n287), .S0(n144), .Y(n189) );
  INVX0_RVT U504 ( .A(a[43]), .Y(n169) );
  MUX21X1_RVT U505 ( .A1(n124), .A2(\u_div/SumTmp[19][23] ), .S0(quotient[19]), 
        .Y(\u_div/PartRem[19][24] ) );
  INVX0_RVT U506 ( .A(\u_div/SumTmp[21][21] ), .Y(n310) );
  MUX21X1_RVT U507 ( .A1(n213), .A2(n311), .S0(quotient[22]), .Y(n236) );
  MUX21X1_RVT U508 ( .A1(n191), .A2(n312), .S0(n109), .Y(n213) );
  INVX0_RVT U509 ( .A(\u_div/SumTmp[23][19] ), .Y(n312) );
  MUX21X1_RVT U510 ( .A1(n170), .A2(n313), .S0(n144), .Y(n191) );
  INVX0_RVT U511 ( .A(\u_div/SumTmp[24][18] ), .Y(n313) );
  INVX0_RVT U512 ( .A(a[42]), .Y(n170) );
  MUX21X1_RVT U513 ( .A1(\u_div/PartRem[19][23] ), .A2(\u_div/SumTmp[18][23] ), 
        .S0(n152), .Y(\u_div/PartRem[18][24] ) );
  MUX21X1_RVT U514 ( .A1(n288), .A2(n337), .S0(quotient[19]), .Y(n336) );
  MUX21X1_RVT U515 ( .A1(n262), .A2(n338), .S0(quotient[20]), .Y(n288) );
  MUX21X1_RVT U516 ( .A1(n237), .A2(n339), .S0(quotient[21]), .Y(n262) );
  INVX0_RVT U517 ( .A(\u_div/SumTmp[21][20] ), .Y(n339) );
  MUX21X1_RVT U518 ( .A1(n214), .A2(n340), .S0(quotient[22]), .Y(n237) );
  INVX0_RVT U519 ( .A(\u_div/SumTmp[22][19] ), .Y(n340) );
  MUX21X1_RVT U520 ( .A1(n192), .A2(n341), .S0(n107), .Y(n214) );
  INVX0_RVT U521 ( .A(\u_div/SumTmp[23][18] ), .Y(n341) );
  MUX21X1_RVT U522 ( .A1(n171), .A2(n342), .S0(n144), .Y(n192) );
  INVX0_RVT U523 ( .A(\u_div/SumTmp[24][17] ), .Y(n342) );
  INVX0_RVT U524 ( .A(a[41]), .Y(n171) );
  MUX21X1_RVT U525 ( .A1(\u_div/PartRem[18][23] ), .A2(\u_div/SumTmp[17][23] ), 
        .S0(n154), .Y(\u_div/PartRem[17][24] ) );
  MUX21X1_RVT U526 ( .A1(n314), .A2(n366), .S0(n152), .Y(n365) );
  MUX21X1_RVT U527 ( .A1(n289), .A2(n367), .S0(quotient[19]), .Y(n314) );
  INVX0_RVT U528 ( .A(\u_div/SumTmp[19][21] ), .Y(n367) );
  MUX21X1_RVT U529 ( .A1(n263), .A2(n368), .S0(quotient[20]), .Y(n289) );
  MUX21X1_RVT U530 ( .A1(n239), .A2(n369), .S0(quotient[21]), .Y(n263) );
  INVX0_RVT U531 ( .A(\u_div/SumTmp[21][19] ), .Y(n369) );
  MUX21X1_RVT U532 ( .A1(n215), .A2(n370), .S0(quotient[22]), .Y(n239) );
  INVX0_RVT U533 ( .A(\u_div/SumTmp[22][18] ), .Y(n370) );
  MUX21X1_RVT U534 ( .A1(n193), .A2(n371), .S0(n106), .Y(n215) );
  INVX0_RVT U535 ( .A(\u_div/SumTmp[23][17] ), .Y(n371) );
  MUX21X1_RVT U536 ( .A1(n172), .A2(n372), .S0(n144), .Y(n193) );
  INVX0_RVT U537 ( .A(\u_div/SumTmp[24][16] ), .Y(n372) );
  INVX0_RVT U538 ( .A(a[40]), .Y(n172) );
  MUX21X1_RVT U539 ( .A1(\u_div/PartRem[17][23] ), .A2(\u_div/SumTmp[16][23] ), 
        .S0(quotient[16]), .Y(\u_div/PartRem[16][24] ) );
  MUX21X1_RVT U540 ( .A1(n343), .A2(n396), .S0(n154), .Y(n395) );
  MUX21X1_RVT U541 ( .A1(n315), .A2(n397), .S0(n152), .Y(n343) );
  INVX0_RVT U542 ( .A(\u_div/SumTmp[18][21] ), .Y(n397) );
  MUX21X1_RVT U543 ( .A1(n290), .A2(n398), .S0(quotient[19]), .Y(n315) );
  INVX0_RVT U544 ( .A(\u_div/SumTmp[19][20] ), .Y(n398) );
  MUX21X1_RVT U545 ( .A1(n265), .A2(n399), .S0(quotient[20]), .Y(n290) );
  INVX0_RVT U546 ( .A(\u_div/SumTmp[20][19] ), .Y(n399) );
  MUX21X1_RVT U547 ( .A1(n240), .A2(n400), .S0(quotient[21]), .Y(n265) );
  INVX0_RVT U548 ( .A(\u_div/SumTmp[21][18] ), .Y(n400) );
  MUX21X1_RVT U549 ( .A1(n216), .A2(n401), .S0(quotient[22]), .Y(n240) );
  INVX0_RVT U550 ( .A(\u_div/SumTmp[22][17] ), .Y(n401) );
  MUX21X1_RVT U551 ( .A1(n194), .A2(n402), .S0(n105), .Y(n216) );
  INVX0_RVT U552 ( .A(\u_div/SumTmp[23][16] ), .Y(n402) );
  MUX21X1_RVT U553 ( .A1(n173), .A2(n403), .S0(n144), .Y(n194) );
  INVX0_RVT U554 ( .A(\u_div/SumTmp[24][15] ), .Y(n403) );
  INVX0_RVT U555 ( .A(a[39]), .Y(n173) );
  MUX21X1_RVT U556 ( .A1(\u_div/PartRem[16][23] ), .A2(\u_div/SumTmp[15][23] ), 
        .S0(n87), .Y(\u_div/PartRem[15][24] ) );
  MUX21X1_RVT U557 ( .A1(n373), .A2(n427), .S0(quotient[16]), .Y(n426) );
  MUX21X1_RVT U558 ( .A1(n344), .A2(n428), .S0(n154), .Y(n373) );
  INVX0_RVT U559 ( .A(\u_div/SumTmp[17][21] ), .Y(n428) );
  MUX21X1_RVT U560 ( .A1(n316), .A2(n429), .S0(n152), .Y(n344) );
  INVX0_RVT U561 ( .A(\u_div/SumTmp[18][20] ), .Y(n429) );
  MUX21X1_RVT U562 ( .A1(n292), .A2(n430), .S0(quotient[19]), .Y(n316) );
  INVX0_RVT U563 ( .A(\u_div/SumTmp[19][19] ), .Y(n430) );
  INVX0_RVT U564 ( .A(\u_div/SumTmp[20][18] ), .Y(n431) );
  MUX21X1_RVT U565 ( .A1(n241), .A2(n432), .S0(quotient[21]), .Y(n266) );
  INVX0_RVT U566 ( .A(\u_div/SumTmp[21][17] ), .Y(n432) );
  MUX21X1_RVT U567 ( .A1(n217), .A2(n433), .S0(quotient[22]), .Y(n241) );
  INVX0_RVT U568 ( .A(\u_div/SumTmp[22][16] ), .Y(n433) );
  MUX21X1_RVT U569 ( .A1(n195), .A2(n434), .S0(n104), .Y(n217) );
  INVX0_RVT U570 ( .A(\u_div/SumTmp[23][15] ), .Y(n434) );
  MUX21X1_RVT U571 ( .A1(n174), .A2(n435), .S0(n144), .Y(n195) );
  INVX0_RVT U572 ( .A(\u_div/SumTmp[24][14] ), .Y(n435) );
  INVX0_RVT U573 ( .A(a[38]), .Y(n174) );
  MUX21X1_RVT U574 ( .A1(n404), .A2(n450), .S0(n87), .Y(n449) );
  INVX0_RVT U575 ( .A(\u_div/SumTmp[15][22] ), .Y(n450) );
  MUX21X1_RVT U576 ( .A1(n374), .A2(n451), .S0(quotient[16]), .Y(n404) );
  INVX0_RVT U577 ( .A(\u_div/SumTmp[16][21] ), .Y(n451) );
  MUX21X1_RVT U578 ( .A1(n345), .A2(n452), .S0(n154), .Y(n374) );
  INVX0_RVT U579 ( .A(\u_div/SumTmp[17][20] ), .Y(n452) );
  MUX21X1_RVT U580 ( .A1(n318), .A2(n453), .S0(n152), .Y(n345) );
  INVX0_RVT U581 ( .A(\u_div/SumTmp[18][19] ), .Y(n453) );
  MUX21X1_RVT U582 ( .A1(n293), .A2(n454), .S0(quotient[19]), .Y(n318) );
  INVX0_RVT U583 ( .A(\u_div/SumTmp[19][18] ), .Y(n454) );
  MUX21X1_RVT U584 ( .A1(n267), .A2(n455), .S0(quotient[20]), .Y(n293) );
  INVX0_RVT U585 ( .A(\u_div/SumTmp[20][17] ), .Y(n455) );
  MUX21X1_RVT U586 ( .A1(n242), .A2(n456), .S0(quotient[21]), .Y(n267) );
  INVX0_RVT U587 ( .A(\u_div/SumTmp[21][16] ), .Y(n456) );
  MUX21X1_RVT U588 ( .A1(n218), .A2(n457), .S0(quotient[22]), .Y(n242) );
  INVX0_RVT U589 ( .A(\u_div/SumTmp[22][15] ), .Y(n457) );
  MUX21X1_RVT U590 ( .A1(n196), .A2(n458), .S0(n103), .Y(n218) );
  INVX0_RVT U591 ( .A(\u_div/SumTmp[23][14] ), .Y(n458) );
  MUX21X1_RVT U592 ( .A1(n175), .A2(n459), .S0(n143), .Y(n196) );
  INVX0_RVT U593 ( .A(\u_div/SumTmp[24][13] ), .Y(n459) );
  INVX0_RVT U594 ( .A(a[37]), .Y(n175) );
  MUX21X1_RVT U595 ( .A1(n405), .A2(n460), .S0(n87), .Y(n436) );
  INVX0_RVT U596 ( .A(\u_div/SumTmp[15][21] ), .Y(n460) );
  MUX21X1_RVT U597 ( .A1(n375), .A2(n461), .S0(quotient[16]), .Y(n405) );
  INVX0_RVT U598 ( .A(\u_div/SumTmp[16][20] ), .Y(n461) );
  MUX21X1_RVT U599 ( .A1(n347), .A2(n462), .S0(n154), .Y(n375) );
  INVX0_RVT U600 ( .A(\u_div/SumTmp[17][19] ), .Y(n462) );
  MUX21X1_RVT U601 ( .A1(n319), .A2(n463), .S0(n152), .Y(n347) );
  INVX0_RVT U602 ( .A(\u_div/SumTmp[18][18] ), .Y(n463) );
  MUX21X1_RVT U603 ( .A1(n294), .A2(n464), .S0(quotient[19]), .Y(n319) );
  INVX0_RVT U604 ( .A(\u_div/SumTmp[19][17] ), .Y(n464) );
  MUX21X1_RVT U605 ( .A1(n268), .A2(n465), .S0(quotient[20]), .Y(n294) );
  MUX21X1_RVT U606 ( .A1(n243), .A2(n466), .S0(quotient[21]), .Y(n268) );
  INVX0_RVT U607 ( .A(\u_div/SumTmp[21][15] ), .Y(n466) );
  MUX21X1_RVT U608 ( .A1(n219), .A2(n467), .S0(quotient[22]), .Y(n243) );
  INVX0_RVT U609 ( .A(\u_div/SumTmp[22][14] ), .Y(n467) );
  MUX21X1_RVT U610 ( .A1(n197), .A2(n468), .S0(quotient[23]), .Y(n219) );
  INVX0_RVT U611 ( .A(\u_div/SumTmp[23][13] ), .Y(n468) );
  MUX21X1_RVT U612 ( .A1(n176), .A2(n469), .S0(n143), .Y(n197) );
  INVX0_RVT U613 ( .A(\u_div/SumTmp[24][12] ), .Y(n469) );
  INVX0_RVT U614 ( .A(a[36]), .Y(n176) );
  MUX21X1_RVT U615 ( .A1(n406), .A2(n470), .S0(n87), .Y(n437) );
  INVX0_RVT U616 ( .A(\u_div/SumTmp[15][20] ), .Y(n470) );
  MUX21X1_RVT U617 ( .A1(n377), .A2(n471), .S0(quotient[16]), .Y(n406) );
  INVX0_RVT U618 ( .A(\u_div/SumTmp[16][19] ), .Y(n471) );
  MUX21X1_RVT U619 ( .A1(n348), .A2(n472), .S0(n154), .Y(n377) );
  MUX21X1_RVT U620 ( .A1(n320), .A2(n473), .S0(n152), .Y(n348) );
  INVX0_RVT U621 ( .A(\u_div/SumTmp[18][17] ), .Y(n473) );
  MUX21X1_RVT U622 ( .A1(n295), .A2(n474), .S0(quotient[19]), .Y(n320) );
  INVX0_RVT U623 ( .A(\u_div/SumTmp[19][16] ), .Y(n474) );
  MUX21X1_RVT U624 ( .A1(n269), .A2(n475), .S0(quotient[20]), .Y(n295) );
  MUX21X1_RVT U625 ( .A1(n244), .A2(n476), .S0(quotient[21]), .Y(n269) );
  INVX0_RVT U626 ( .A(\u_div/SumTmp[21][14] ), .Y(n476) );
  MUX21X1_RVT U627 ( .A1(n220), .A2(n477), .S0(n146), .Y(n244) );
  INVX0_RVT U628 ( .A(\u_div/SumTmp[22][13] ), .Y(n477) );
  MUX21X1_RVT U629 ( .A1(n198), .A2(n478), .S0(n114), .Y(n220) );
  INVX0_RVT U630 ( .A(\u_div/SumTmp[23][12] ), .Y(n478) );
  MUX21X1_RVT U631 ( .A1(n177), .A2(n479), .S0(n143), .Y(n198) );
  INVX0_RVT U632 ( .A(\u_div/SumTmp[24][11] ), .Y(n479) );
  INVX0_RVT U633 ( .A(a[35]), .Y(n177) );
  MUX21X1_RVT U634 ( .A1(n408), .A2(n480), .S0(n87), .Y(n438) );
  INVX0_RVT U635 ( .A(\u_div/SumTmp[15][19] ), .Y(n480) );
  MUX21X1_RVT U636 ( .A1(n349), .A2(n482), .S0(n154), .Y(n378) );
  INVX0_RVT U637 ( .A(\u_div/SumTmp[17][17] ), .Y(n482) );
  MUX21X1_RVT U638 ( .A1(n321), .A2(n483), .S0(n152), .Y(n349) );
  INVX0_RVT U639 ( .A(\u_div/SumTmp[18][16] ), .Y(n483) );
  MUX21X1_RVT U640 ( .A1(n296), .A2(n484), .S0(quotient[19]), .Y(n321) );
  INVX0_RVT U641 ( .A(\u_div/SumTmp[19][15] ), .Y(n484) );
  MUX21X1_RVT U642 ( .A1(n270), .A2(n485), .S0(quotient[20]), .Y(n296) );
  INVX0_RVT U643 ( .A(\u_div/SumTmp[20][14] ), .Y(n485) );
  MUX21X1_RVT U644 ( .A1(n245), .A2(n486), .S0(quotient[21]), .Y(n270) );
  INVX0_RVT U645 ( .A(\u_div/SumTmp[21][13] ), .Y(n486) );
  INVX0_RVT U646 ( .A(\u_div/SumTmp[22][12] ), .Y(n487) );
  MUX21X1_RVT U647 ( .A1(n199), .A2(n488), .S0(quotient[23]), .Y(n221) );
  INVX0_RVT U648 ( .A(\u_div/SumTmp[23][11] ), .Y(n488) );
  MUX21X1_RVT U649 ( .A1(n178), .A2(n489), .S0(n143), .Y(n199) );
  INVX0_RVT U650 ( .A(\u_div/SumTmp[24][10] ), .Y(n489) );
  INVX0_RVT U651 ( .A(a[34]), .Y(n178) );
  MUX21X1_RVT U652 ( .A1(n393), .A2(n490), .S0(n87), .Y(n423) );
  INVX0_RVT U653 ( .A(\u_div/SumTmp[15][3] ), .Y(n490) );
  MUX21X1_RVT U654 ( .A1(n364), .A2(n491), .S0(quotient[16]), .Y(n393) );
  INVX0_RVT U655 ( .A(\u_div/SumTmp[16][2] ), .Y(n491) );
  MUX21X1_RVT U656 ( .A1(n346), .A2(n492), .S0(n154), .Y(n364) );
  INVX0_RVT U657 ( .A(\u_div/SumTmp[17][1] ), .Y(n492) );
  MUX21X1_RVT U658 ( .A1(n394), .A2(n493), .S0(n87), .Y(n424) );
  INVX0_RVT U659 ( .A(\u_div/SumTmp[15][2] ), .Y(n493) );
  MUX21X1_RVT U660 ( .A1(n376), .A2(n494), .S0(quotient[16]), .Y(n394) );
  INVX0_RVT U661 ( .A(\u_div/SumTmp[16][1] ), .Y(n494) );
  MUX21X1_RVT U662 ( .A1(n407), .A2(n495), .S0(n87), .Y(n425) );
  INVX0_RVT U663 ( .A(\u_div/SumTmp[15][1] ), .Y(n495) );
  MUX21X1_RVT U664 ( .A1(n409), .A2(n496), .S0(n87), .Y(n439) );
  INVX0_RVT U665 ( .A(\u_div/SumTmp[15][18] ), .Y(n496) );
  MUX21X1_RVT U666 ( .A1(n379), .A2(n497), .S0(quotient[16]), .Y(n409) );
  INVX0_RVT U667 ( .A(\u_div/SumTmp[16][17] ), .Y(n497) );
  MUX21X1_RVT U668 ( .A1(n350), .A2(n498), .S0(n154), .Y(n379) );
  INVX0_RVT U669 ( .A(\u_div/SumTmp[17][16] ), .Y(n498) );
  MUX21X1_RVT U670 ( .A1(n322), .A2(n499), .S0(n152), .Y(n350) );
  INVX0_RVT U671 ( .A(\u_div/SumTmp[18][15] ), .Y(n499) );
  MUX21X1_RVT U672 ( .A1(n297), .A2(n500), .S0(quotient[19]), .Y(n322) );
  INVX0_RVT U673 ( .A(\u_div/SumTmp[19][14] ), .Y(n500) );
  MUX21X1_RVT U674 ( .A1(n271), .A2(n501), .S0(n148), .Y(n297) );
  INVX0_RVT U675 ( .A(\u_div/SumTmp[20][13] ), .Y(n501) );
  MUX21X1_RVT U676 ( .A1(n246), .A2(n502), .S0(quotient[21]), .Y(n271) );
  INVX0_RVT U677 ( .A(\u_div/SumTmp[21][12] ), .Y(n502) );
  INVX0_RVT U678 ( .A(\u_div/SumTmp[22][11] ), .Y(n503) );
  MUX21X1_RVT U679 ( .A1(n200), .A2(n504), .S0(quotient[23]), .Y(n222) );
  INVX0_RVT U680 ( .A(\u_div/SumTmp[23][10] ), .Y(n504) );
  MUX21X1_RVT U681 ( .A1(n157), .A2(n505), .S0(n143), .Y(n200) );
  INVX0_RVT U682 ( .A(\u_div/SumTmp[24][9] ), .Y(n505) );
  INVX0_RVT U683 ( .A(a[33]), .Y(n157) );
  MUX21X1_RVT U684 ( .A1(n410), .A2(n506), .S0(n87), .Y(n440) );
  INVX0_RVT U685 ( .A(\u_div/SumTmp[15][17] ), .Y(n506) );
  MUX21X1_RVT U686 ( .A1(n380), .A2(n507), .S0(quotient[16]), .Y(n410) );
  INVX0_RVT U687 ( .A(\u_div/SumTmp[16][16] ), .Y(n507) );
  MUX21X1_RVT U688 ( .A1(n351), .A2(n508), .S0(n154), .Y(n380) );
  INVX0_RVT U689 ( .A(\u_div/SumTmp[17][15] ), .Y(n508) );
  MUX21X1_RVT U690 ( .A1(n323), .A2(n509), .S0(n152), .Y(n351) );
  INVX0_RVT U691 ( .A(\u_div/SumTmp[18][14] ), .Y(n509) );
  MUX21X1_RVT U692 ( .A1(n298), .A2(n510), .S0(n100), .Y(n323) );
  INVX0_RVT U693 ( .A(\u_div/SumTmp[19][13] ), .Y(n510) );
  MUX21X1_RVT U694 ( .A1(n272), .A2(n511), .S0(n148), .Y(n298) );
  INVX0_RVT U695 ( .A(\u_div/SumTmp[20][12] ), .Y(n511) );
  MUX21X1_RVT U696 ( .A1(n247), .A2(n512), .S0(quotient[21]), .Y(n272) );
  INVX0_RVT U697 ( .A(\u_div/SumTmp[21][11] ), .Y(n512) );
  INVX0_RVT U698 ( .A(\u_div/SumTmp[22][10] ), .Y(n513) );
  MUX21X1_RVT U699 ( .A1(n179), .A2(n514), .S0(quotient[23]), .Y(n223) );
  INVX0_RVT U700 ( .A(\u_div/SumTmp[23][9] ), .Y(n514) );
  MUX21X1_RVT U701 ( .A1(n158), .A2(n515), .S0(n143), .Y(n179) );
  INVX0_RVT U702 ( .A(\u_div/SumTmp[24][8] ), .Y(n515) );
  INVX0_RVT U703 ( .A(a[32]), .Y(n158) );
  MUX21X1_RVT U704 ( .A1(n411), .A2(n516), .S0(n87), .Y(n441) );
  INVX0_RVT U705 ( .A(\u_div/SumTmp[15][16] ), .Y(n516) );
  MUX21X1_RVT U706 ( .A1(n381), .A2(n517), .S0(quotient[16]), .Y(n411) );
  INVX0_RVT U707 ( .A(\u_div/SumTmp[16][15] ), .Y(n517) );
  MUX21X1_RVT U708 ( .A1(n352), .A2(n518), .S0(n154), .Y(n381) );
  INVX0_RVT U709 ( .A(\u_div/SumTmp[17][14] ), .Y(n518) );
  MUX21X1_RVT U710 ( .A1(n324), .A2(n519), .S0(n152), .Y(n352) );
  INVX0_RVT U711 ( .A(\u_div/SumTmp[18][13] ), .Y(n519) );
  MUX21X1_RVT U712 ( .A1(n299), .A2(n520), .S0(n100), .Y(n324) );
  INVX0_RVT U713 ( .A(\u_div/SumTmp[19][12] ), .Y(n520) );
  MUX21X1_RVT U714 ( .A1(n273), .A2(n521), .S0(n148), .Y(n299) );
  INVX0_RVT U715 ( .A(\u_div/SumTmp[20][11] ), .Y(n521) );
  MUX21X1_RVT U716 ( .A1(n248), .A2(n522), .S0(quotient[21]), .Y(n273) );
  INVX0_RVT U717 ( .A(\u_div/SumTmp[21][10] ), .Y(n522) );
  INVX0_RVT U718 ( .A(\u_div/SumTmp[22][9] ), .Y(n523) );
  MUX21X1_RVT U719 ( .A1(n180), .A2(n524), .S0(n114), .Y(n201) );
  INVX0_RVT U720 ( .A(\u_div/SumTmp[23][8] ), .Y(n524) );
  MUX21X1_RVT U721 ( .A1(n159), .A2(n525), .S0(n143), .Y(n180) );
  INVX0_RVT U722 ( .A(\u_div/SumTmp[24][7] ), .Y(n525) );
  INVX0_RVT U723 ( .A(a[31]), .Y(n159) );
  MUX21X1_RVT U724 ( .A1(n412), .A2(n526), .S0(n87), .Y(n442) );
  INVX0_RVT U725 ( .A(\u_div/SumTmp[15][15] ), .Y(n526) );
  MUX21X1_RVT U726 ( .A1(n382), .A2(n527), .S0(quotient[16]), .Y(n412) );
  INVX0_RVT U727 ( .A(\u_div/SumTmp[16][14] ), .Y(n527) );
  MUX21X1_RVT U728 ( .A1(n353), .A2(n528), .S0(n154), .Y(n382) );
  INVX0_RVT U729 ( .A(\u_div/SumTmp[17][13] ), .Y(n528) );
  MUX21X1_RVT U730 ( .A1(n325), .A2(n529), .S0(n152), .Y(n353) );
  MUX21X1_RVT U731 ( .A1(n300), .A2(n530), .S0(n100), .Y(n325) );
  INVX0_RVT U732 ( .A(\u_div/SumTmp[19][11] ), .Y(n530) );
  MUX21X1_RVT U733 ( .A1(n274), .A2(n531), .S0(n148), .Y(n300) );
  INVX0_RVT U734 ( .A(\u_div/SumTmp[20][10] ), .Y(n531) );
  MUX21X1_RVT U735 ( .A1(n224), .A2(n532), .S0(quotient[21]), .Y(n274) );
  INVX0_RVT U736 ( .A(\u_div/SumTmp[21][9] ), .Y(n532) );
  INVX0_RVT U737 ( .A(\u_div/SumTmp[22][8] ), .Y(n533) );
  MUX21X1_RVT U738 ( .A1(n181), .A2(n534), .S0(n112), .Y(n202) );
  INVX0_RVT U739 ( .A(\u_div/SumTmp[23][7] ), .Y(n534) );
  MUX21X1_RVT U740 ( .A1(n160), .A2(n535), .S0(n143), .Y(n181) );
  INVX0_RVT U741 ( .A(\u_div/SumTmp[24][6] ), .Y(n535) );
  INVX0_RVT U742 ( .A(a[30]), .Y(n160) );
  MUX21X1_RVT U743 ( .A1(n413), .A2(n536), .S0(quotient[15]), .Y(n443) );
  MUX21X1_RVT U744 ( .A1(n383), .A2(n537), .S0(quotient[16]), .Y(n413) );
  INVX0_RVT U745 ( .A(\u_div/SumTmp[16][13] ), .Y(n537) );
  MUX21X1_RVT U746 ( .A1(n354), .A2(n538), .S0(quotient[17]), .Y(n383) );
  INVX0_RVT U747 ( .A(\u_div/SumTmp[17][12] ), .Y(n538) );
  MUX21X1_RVT U748 ( .A1(n326), .A2(n539), .S0(quotient[18]), .Y(n354) );
  INVX0_RVT U749 ( .A(\u_div/SumTmp[18][11] ), .Y(n539) );
  MUX21X1_RVT U750 ( .A1(n301), .A2(n43), .S0(n100), .Y(n326) );
  MUX21X1_RVT U751 ( .A1(n249), .A2(n540), .S0(n148), .Y(n301) );
  MUX21X1_RVT U752 ( .A1(n225), .A2(n541), .S0(quotient[21]), .Y(n249) );
  INVX0_RVT U753 ( .A(\u_div/SumTmp[21][8] ), .Y(n541) );
  INVX0_RVT U754 ( .A(\u_div/SumTmp[22][7] ), .Y(n542) );
  MUX21X1_RVT U755 ( .A1(n182), .A2(n543), .S0(n111), .Y(n203) );
  INVX0_RVT U756 ( .A(\u_div/SumTmp[23][6] ), .Y(n543) );
  MUX21X1_RVT U757 ( .A1(n161), .A2(n544), .S0(n143), .Y(n182) );
  INVX0_RVT U758 ( .A(\u_div/SumTmp[24][5] ), .Y(n544) );
  INVX0_RVT U759 ( .A(a[29]), .Y(n161) );
  MUX21X1_RVT U760 ( .A1(n414), .A2(n545), .S0(quotient[15]), .Y(n444) );
  INVX0_RVT U761 ( .A(\u_div/SumTmp[15][13] ), .Y(n545) );
  MUX21X1_RVT U762 ( .A1(n384), .A2(n546), .S0(quotient[16]), .Y(n414) );
  INVX0_RVT U763 ( .A(\u_div/SumTmp[16][12] ), .Y(n546) );
  MUX21X1_RVT U764 ( .A1(n355), .A2(n547), .S0(quotient[17]), .Y(n384) );
  INVX0_RVT U765 ( .A(\u_div/SumTmp[17][11] ), .Y(n547) );
  MUX21X1_RVT U766 ( .A1(n327), .A2(n548), .S0(quotient[18]), .Y(n355) );
  INVX0_RVT U767 ( .A(\u_div/SumTmp[18][10] ), .Y(n548) );
  MUX21X1_RVT U768 ( .A1(n275), .A2(n549), .S0(n100), .Y(n327) );
  INVX0_RVT U769 ( .A(\u_div/SumTmp[19][9] ), .Y(n549) );
  MUX21X1_RVT U770 ( .A1(n250), .A2(n550), .S0(n148), .Y(n275) );
  INVX0_RVT U771 ( .A(\u_div/SumTmp[20][8] ), .Y(n550) );
  MUX21X1_RVT U772 ( .A1(n226), .A2(n551), .S0(quotient[21]), .Y(n250) );
  INVX0_RVT U773 ( .A(\u_div/SumTmp[21][7] ), .Y(n551) );
  INVX0_RVT U774 ( .A(\u_div/SumTmp[22][6] ), .Y(n552) );
  MUX21X1_RVT U775 ( .A1(n183), .A2(n553), .S0(n110), .Y(n204) );
  INVX0_RVT U776 ( .A(\u_div/SumTmp[23][5] ), .Y(n553) );
  MUX21X1_RVT U777 ( .A1(n162), .A2(n554), .S0(n143), .Y(n183) );
  INVX0_RVT U778 ( .A(\u_div/SumTmp[24][4] ), .Y(n554) );
  INVX0_RVT U779 ( .A(a[28]), .Y(n162) );
  MUX21X1_RVT U780 ( .A1(n415), .A2(n555), .S0(quotient[15]), .Y(n445) );
  MUX21X1_RVT U781 ( .A1(n385), .A2(n556), .S0(quotient[16]), .Y(n415) );
  INVX0_RVT U782 ( .A(\u_div/SumTmp[16][11] ), .Y(n556) );
  MUX21X1_RVT U783 ( .A1(n356), .A2(n557), .S0(quotient[17]), .Y(n385) );
  INVX0_RVT U784 ( .A(\u_div/SumTmp[17][10] ), .Y(n557) );
  MUX21X1_RVT U785 ( .A1(n302), .A2(n558), .S0(quotient[18]), .Y(n356) );
  INVX0_RVT U786 ( .A(\u_div/SumTmp[18][9] ), .Y(n558) );
  MUX21X1_RVT U787 ( .A1(n276), .A2(n559), .S0(n100), .Y(n302) );
  INVX0_RVT U788 ( .A(\u_div/SumTmp[19][8] ), .Y(n559) );
  MUX21X1_RVT U789 ( .A1(n251), .A2(n560), .S0(n148), .Y(n276) );
  INVX0_RVT U790 ( .A(\u_div/SumTmp[20][7] ), .Y(n560) );
  MUX21X1_RVT U791 ( .A1(n227), .A2(n561), .S0(quotient[21]), .Y(n251) );
  INVX0_RVT U792 ( .A(\u_div/SumTmp[21][6] ), .Y(n561) );
  INVX0_RVT U793 ( .A(\u_div/SumTmp[22][5] ), .Y(n562) );
  MUX21X1_RVT U794 ( .A1(n184), .A2(n563), .S0(n109), .Y(n205) );
  INVX0_RVT U795 ( .A(\u_div/SumTmp[23][4] ), .Y(n563) );
  MUX21X1_RVT U796 ( .A1(n163), .A2(n564), .S0(n143), .Y(n184) );
  INVX0_RVT U797 ( .A(\u_div/SumTmp[24][3] ), .Y(n564) );
  INVX0_RVT U798 ( .A(a[27]), .Y(n163) );
  MUX21X1_RVT U799 ( .A1(n416), .A2(n565), .S0(quotient[15]), .Y(n446) );
  INVX0_RVT U800 ( .A(\u_div/SumTmp[15][11] ), .Y(n565) );
  MUX21X1_RVT U801 ( .A1(n386), .A2(n566), .S0(quotient[16]), .Y(n416) );
  INVX0_RVT U802 ( .A(\u_div/SumTmp[16][10] ), .Y(n566) );
  MUX21X1_RVT U803 ( .A1(n328), .A2(n567), .S0(quotient[17]), .Y(n386) );
  INVX0_RVT U804 ( .A(\u_div/SumTmp[17][9] ), .Y(n567) );
  MUX21X1_RVT U805 ( .A1(n303), .A2(n568), .S0(quotient[18]), .Y(n328) );
  INVX0_RVT U806 ( .A(\u_div/SumTmp[18][8] ), .Y(n568) );
  MUX21X1_RVT U807 ( .A1(n277), .A2(n569), .S0(n100), .Y(n303) );
  INVX0_RVT U808 ( .A(\u_div/SumTmp[19][7] ), .Y(n569) );
  MUX21X1_RVT U809 ( .A1(n252), .A2(n570), .S0(n148), .Y(n277) );
  INVX0_RVT U810 ( .A(\u_div/SumTmp[20][6] ), .Y(n570) );
  MUX21X1_RVT U811 ( .A1(n228), .A2(n571), .S0(quotient[21]), .Y(n252) );
  INVX0_RVT U812 ( .A(\u_div/SumTmp[21][5] ), .Y(n571) );
  INVX0_RVT U813 ( .A(\u_div/SumTmp[22][4] ), .Y(n572) );
  MUX21X1_RVT U814 ( .A1(n185), .A2(n573), .S0(n107), .Y(n206) );
  INVX0_RVT U815 ( .A(\u_div/SumTmp[23][3] ), .Y(n573) );
  MUX21X1_RVT U816 ( .A1(n164), .A2(n574), .S0(n143), .Y(n185) );
  INVX0_RVT U817 ( .A(\u_div/SumTmp[24][2] ), .Y(n574) );
  INVX0_RVT U818 ( .A(a[26]), .Y(n164) );
  MUX21X1_RVT U819 ( .A1(n417), .A2(n575), .S0(quotient[15]), .Y(n447) );
  INVX0_RVT U820 ( .A(\u_div/SumTmp[15][10] ), .Y(n575) );
  MUX21X1_RVT U821 ( .A1(n357), .A2(n576), .S0(quotient[16]), .Y(n417) );
  INVX0_RVT U822 ( .A(\u_div/SumTmp[16][9] ), .Y(n576) );
  MUX21X1_RVT U823 ( .A1(n329), .A2(n577), .S0(quotient[17]), .Y(n357) );
  INVX0_RVT U824 ( .A(\u_div/SumTmp[17][8] ), .Y(n577) );
  MUX21X1_RVT U825 ( .A1(n304), .A2(n578), .S0(quotient[18]), .Y(n329) );
  INVX0_RVT U826 ( .A(\u_div/SumTmp[18][7] ), .Y(n578) );
  MUX21X1_RVT U827 ( .A1(n278), .A2(n579), .S0(n100), .Y(n304) );
  INVX0_RVT U828 ( .A(\u_div/SumTmp[19][6] ), .Y(n579) );
  MUX21X1_RVT U829 ( .A1(n253), .A2(n580), .S0(n148), .Y(n278) );
  INVX0_RVT U830 ( .A(\u_div/SumTmp[20][5] ), .Y(n580) );
  MUX21X1_RVT U831 ( .A1(n229), .A2(n581), .S0(quotient[21]), .Y(n253) );
  INVX0_RVT U832 ( .A(\u_div/SumTmp[21][4] ), .Y(n581) );
  INVX0_RVT U833 ( .A(\u_div/SumTmp[22][3] ), .Y(n582) );
  MUX21X1_RVT U834 ( .A1(n186), .A2(n583), .S0(n106), .Y(n207) );
  INVX0_RVT U835 ( .A(\u_div/SumTmp[23][2] ), .Y(n583) );
  MUX21X1_RVT U836 ( .A1(n168), .A2(n584), .S0(n143), .Y(n186) );
  INVX0_RVT U837 ( .A(a[25]), .Y(n168) );
  MUX21X1_RVT U838 ( .A1(n387), .A2(n585), .S0(quotient[15]), .Y(n448) );
  INVX0_RVT U839 ( .A(\u_div/SumTmp[15][9] ), .Y(n585) );
  MUX21X1_RVT U840 ( .A1(n358), .A2(n586), .S0(quotient[16]), .Y(n387) );
  INVX0_RVT U841 ( .A(\u_div/SumTmp[16][8] ), .Y(n586) );
  MUX21X1_RVT U842 ( .A1(n330), .A2(n587), .S0(quotient[17]), .Y(n358) );
  INVX0_RVT U843 ( .A(\u_div/SumTmp[17][7] ), .Y(n587) );
  MUX21X1_RVT U844 ( .A1(n305), .A2(n588), .S0(quotient[18]), .Y(n330) );
  INVX0_RVT U845 ( .A(\u_div/SumTmp[18][6] ), .Y(n588) );
  MUX21X1_RVT U846 ( .A1(n279), .A2(n589), .S0(n100), .Y(n305) );
  INVX0_RVT U847 ( .A(\u_div/SumTmp[19][5] ), .Y(n589) );
  MUX21X1_RVT U848 ( .A1(n254), .A2(n590), .S0(n148), .Y(n279) );
  INVX0_RVT U849 ( .A(\u_div/SumTmp[20][4] ), .Y(n590) );
  MUX21X1_RVT U850 ( .A1(n230), .A2(n591), .S0(quotient[21]), .Y(n254) );
  INVX0_RVT U851 ( .A(\u_div/SumTmp[21][3] ), .Y(n591) );
  INVX0_RVT U852 ( .A(\u_div/SumTmp[22][2] ), .Y(n592) );
  MUX21X1_RVT U853 ( .A1(n190), .A2(n593), .S0(n105), .Y(n208) );
  INVX0_RVT U854 ( .A(\u_div/SumTmp[23][1] ), .Y(n593) );
  MUX21X2_RVT U855 ( .A1(n594), .A2(n125), .S0(n143), .Y(n190) );
  MUX21X1_RVT U856 ( .A1(n388), .A2(n595), .S0(quotient[15]), .Y(n418) );
  INVX0_RVT U857 ( .A(\u_div/SumTmp[15][8] ), .Y(n595) );
  MUX21X1_RVT U858 ( .A1(n359), .A2(n596), .S0(quotient[16]), .Y(n388) );
  INVX0_RVT U859 ( .A(\u_div/SumTmp[16][7] ), .Y(n596) );
  MUX21X1_RVT U860 ( .A1(n331), .A2(n597), .S0(quotient[17]), .Y(n359) );
  INVX0_RVT U861 ( .A(\u_div/SumTmp[17][6] ), .Y(n597) );
  MUX21X1_RVT U862 ( .A1(n306), .A2(n598), .S0(quotient[18]), .Y(n331) );
  INVX0_RVT U863 ( .A(\u_div/SumTmp[18][5] ), .Y(n598) );
  MUX21X1_RVT U864 ( .A1(n280), .A2(n599), .S0(n100), .Y(n306) );
  INVX0_RVT U865 ( .A(\u_div/SumTmp[19][4] ), .Y(n599) );
  MUX21X1_RVT U866 ( .A1(n255), .A2(n600), .S0(n148), .Y(n280) );
  MUX21X1_RVT U867 ( .A1(n231), .A2(n601), .S0(quotient[21]), .Y(n255) );
  INVX0_RVT U868 ( .A(\u_div/SumTmp[21][2] ), .Y(n601) );
  INVX0_RVT U869 ( .A(\u_div/SumTmp[23][0] ), .Y(n602) );
  MUX21X1_RVT U870 ( .A1(n389), .A2(n603), .S0(quotient[15]), .Y(n419) );
  INVX0_RVT U871 ( .A(\u_div/SumTmp[15][7] ), .Y(n603) );
  MUX21X1_RVT U872 ( .A1(n360), .A2(n604), .S0(quotient[16]), .Y(n389) );
  INVX0_RVT U873 ( .A(\u_div/SumTmp[16][6] ), .Y(n604) );
  MUX21X1_RVT U874 ( .A1(n332), .A2(n605), .S0(quotient[17]), .Y(n360) );
  INVX0_RVT U875 ( .A(\u_div/SumTmp[17][5] ), .Y(n605) );
  MUX21X1_RVT U876 ( .A1(n307), .A2(n606), .S0(quotient[18]), .Y(n332) );
  INVX0_RVT U877 ( .A(\u_div/SumTmp[18][4] ), .Y(n606) );
  MUX21X1_RVT U878 ( .A1(n281), .A2(n607), .S0(n100), .Y(n307) );
  INVX0_RVT U879 ( .A(\u_div/SumTmp[19][3] ), .Y(n607) );
  MUX21X1_RVT U880 ( .A1(n256), .A2(n608), .S0(n148), .Y(n281) );
  MUX21X1_RVT U881 ( .A1(n68), .A2(n609), .S0(quotient[21]), .Y(n256) );
  INVX0_RVT U882 ( .A(\u_div/SumTmp[21][1] ), .Y(n609) );
  INVX0_RVT U883 ( .A(\u_div/SumTmp[22][0] ), .Y(n610) );
  MUX21X1_RVT U884 ( .A1(n390), .A2(n611), .S0(quotient[15]), .Y(n420) );
  INVX0_RVT U885 ( .A(\u_div/SumTmp[15][6] ), .Y(n611) );
  MUX21X1_RVT U886 ( .A1(n361), .A2(n612), .S0(quotient[16]), .Y(n390) );
  INVX0_RVT U887 ( .A(\u_div/SumTmp[16][5] ), .Y(n612) );
  MUX21X1_RVT U888 ( .A1(n333), .A2(n613), .S0(quotient[17]), .Y(n361) );
  INVX0_RVT U889 ( .A(\u_div/SumTmp[17][4] ), .Y(n613) );
  MUX21X1_RVT U890 ( .A1(n308), .A2(n614), .S0(quotient[18]), .Y(n333) );
  INVX0_RVT U891 ( .A(\u_div/SumTmp[18][3] ), .Y(n614) );
  MUX21X1_RVT U892 ( .A1(n282), .A2(n615), .S0(n100), .Y(n308) );
  INVX0_RVT U893 ( .A(\u_div/SumTmp[19][2] ), .Y(n615) );
  MUX21X1_RVT U894 ( .A1(n264), .A2(n616), .S0(n148), .Y(n282) );
  INVX0_RVT U895 ( .A(\u_div/SumTmp[20][1] ), .Y(n616) );
  INVX0_RVT U896 ( .A(\u_div/SumTmp[21][0] ), .Y(n617) );
  MUX21X1_RVT U897 ( .A1(n391), .A2(n618), .S0(quotient[15]), .Y(n421) );
  INVX0_RVT U898 ( .A(\u_div/SumTmp[15][5] ), .Y(n618) );
  MUX21X1_RVT U899 ( .A1(n362), .A2(n619), .S0(quotient[16]), .Y(n391) );
  INVX0_RVT U900 ( .A(\u_div/SumTmp[16][4] ), .Y(n619) );
  MUX21X1_RVT U901 ( .A1(n334), .A2(n620), .S0(quotient[17]), .Y(n362) );
  INVX0_RVT U902 ( .A(\u_div/SumTmp[17][3] ), .Y(n620) );
  MUX21X1_RVT U903 ( .A1(n291), .A2(n622), .S0(n100), .Y(n309) );
  INVX0_RVT U904 ( .A(\u_div/SumTmp[19][1] ), .Y(n622) );
  INVX0_RVT U905 ( .A(\u_div/SumTmp[20][0] ), .Y(n623) );
  MUX21X1_RVT U906 ( .A1(n392), .A2(n624), .S0(n87), .Y(n422) );
  INVX0_RVT U907 ( .A(\u_div/SumTmp[15][4] ), .Y(n624) );
  MUX21X1_RVT U908 ( .A1(n363), .A2(n625), .S0(quotient[16]), .Y(n392) );
  INVX0_RVT U909 ( .A(\u_div/SumTmp[16][3] ), .Y(n625) );
  MUX21X1_RVT U910 ( .A1(n335), .A2(n626), .S0(n154), .Y(n363) );
  INVX0_RVT U911 ( .A(\u_div/SumTmp[17][2] ), .Y(n626) );
  MUX21X1_RVT U912 ( .A1(n317), .A2(n627), .S0(n152), .Y(n335) );
  INVX0_RVT U913 ( .A(\u_div/SumTmp[18][1] ), .Y(n627) );
  INVX0_RVT U914 ( .A(\u_div/SumTmp[19][0] ), .Y(n628) );
endmodule


module FPU_CAL ( clk, start, A, B, sel, round_mode, error, over_flow, Y );
  input [31:0] A;
  input [31:0] B;
  input [1:0] sel;
  output [31:0] Y;
  input clk, start, round_mode;
  output error, over_flow;
  wire   N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123,
         N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134,
         N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153,
         N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164,
         N165, N166, N167, N172, N173, N174, N175, N176, N177, N178, N179,
         N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190,
         N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201,
         N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212,
         N213, N214, N215, N216, N217, N218, N219, N220, N221, N248, N249,
         N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260,
         N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271,
         N272, N330, N331, N332, N333, N334, N335, N336, N337, N338, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374,
         N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385,
         N386, N387, N388, N389, N390, N391, N392, N393, N394, N395, N396,
         N397, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N418, N419, N420, N421, N422, N423, N424, N438, N439, N440,
         N441, N442, N443, N444, N445, N446, N493, N494, N495, N496, N497,
         N498, N499, N500, N501, N505, N506, N507, N508, N509, N510, N511,
         N512, N513, N516, N519, N520, N521, N522, N523, N524, N525, N526,
         N527, N536, N545, N573, N574, N575, N576, N577, N578, N579, N580,
         N604, N605, N606, N607, N608, N609, N610, N611, N634, N635, N636,
         N637, N638, N639, N640, N641, n140, n141, n143, n202, n211, n214,
         n217, n220, n223, n226, n323, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n500, n501, n503, n504, n505, n506, n507, n509, n510, n511,
         n512, n514, n515, n516, n517, n518, n520, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, N350, N349, N348, N347,
         N346, N345, N344, N437, N492, N491, N490, N489, N488, N487, N486,
         N485, N484, \sub_143/carry[2] , \sub_143/carry[3] ,
         \sub_143/carry[4] , \sub_143/carry[5] , \sub_143/carry[6] ,
         \sub_143/carry[7] , \sub_1_root_sub_0_root_sub_122/carry[2] ,
         \sub_1_root_sub_0_root_sub_122/carry[3] ,
         \sub_1_root_sub_0_root_sub_122/carry[4] ,
         \sub_1_root_sub_0_root_sub_122/carry[5] ,
         \sub_1_root_sub_0_root_sub_122/carry[6] ,
         \sub_1_root_sub_0_root_sub_122/carry[7] ,
         \sub_1_root_add_170/carry[8] , \sub_1_root_add_170/carry[7] ,
         \sub_1_root_add_170/carry[5] , \sub_1_root_add_170/carry[4] ,
         \sub_1_root_add_170/carry[3] , \sub_1_root_add_170/carry[2] ,
         \sub_1_root_add_170/carry[1] , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n122, n124, n126, n128, n130, n132, n134,
         n136, n137, n138, n139, n142, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n203, n204, n205,
         n206, n207, n208, n209, n210, n212, n213, n215, n216, n218, n219,
         n221, n222, n224, n225, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n499, n502, n508, n513, n519, n521, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752;
  wire   [24:0] M_sum;
  wire   [22:0] result;
  wire   [4:0] shifted;
  wire   [2:0] next_state;
  wire   [8:0] E;
  wire   [47:0] M1M2;
  wire   [47:0] div;
  wire   [23:0] divider;
  wire   [23:15] quotient;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52;
  assign Y[14] = 1'b0;
  assign Y[13] = 1'b0;
  assign Y[12] = 1'b0;
  assign Y[11] = 1'b0;
  assign Y[10] = 1'b0;
  assign Y[9] = 1'b0;
  assign Y[8] = 1'b0;
  assign Y[7] = 1'b0;
  assign Y[6] = 1'b0;
  assign Y[5] = 1'b0;
  assign Y[4] = 1'b0;
  assign Y[3] = 1'b0;
  assign Y[2] = 1'b0;
  assign Y[1] = 1'b0;
  assign Y[0] = 1'b0;
  assign N437 = B[30];

  DFFSSRX1_RVT \E_reg[8]  ( .D(n323), .SETB(n745), .RSTB(1'b1), .CLK(clk), .Q(
        n285), .QN(n741) );
  DFFSSRX1_RVT \Y_reg[21]  ( .D(n202), .SETB(n746), .RSTB(1'b1), .CLK(clk), 
        .Q(Y[21]) );
  DFFSSRX1_RVT \Y_reg[20]  ( .D(n211), .SETB(n747), .RSTB(1'b1), .CLK(clk), 
        .Q(Y[20]) );
  DFFSSRX1_RVT \Y_reg[19]  ( .D(n214), .SETB(n748), .RSTB(1'b1), .CLK(clk), 
        .Q(Y[19]) );
  DFFSSRX1_RVT \Y_reg[18]  ( .D(n217), .SETB(n749), .RSTB(1'b1), .CLK(clk), 
        .Q(Y[18]) );
  DFFSSRX1_RVT \Y_reg[17]  ( .D(n220), .SETB(n750), .RSTB(1'b1), .CLK(clk), 
        .Q(Y[17]) );
  DFFSSRX1_RVT \Y_reg[16]  ( .D(n223), .SETB(n751), .RSTB(1'b1), .CLK(clk), 
        .Q(Y[16]) );
  DFFSSRX1_RVT \Y_reg[15]  ( .D(n226), .SETB(n752), .RSTB(1'b1), .CLK(clk), 
        .Q(Y[15]) );
  FPU_normalize fpu_normalize ( .src({n229, n231, n233, n235, n237, n239, n241, 
        n243, n245, M_sum[15], n288, n247, n249, n251, n252, n254, M_sum[8], 
        n255, n256, n258, n260, n262, n264, n266, n268}), .result({
        result[22:15], SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14}), .shifted(shifted) );
  FPU_CAL_DW01_inc_0 add_232 ( .A(quotient[23:16]), .SUM({N641, N640, N639, 
        N638, N637, N636, N635, N634}) );
  FPU_CAL_DW01_inc_1 add_218 ( .A(M1M2[46:39]), .SUM({N611, N610, N609, N608, 
        N607, N606, N605, N604}) );
  FPU_CAL_DW01_inc_2 add_204 ( .A(result[22:15]), .SUM({N580, N579, N578, N577, 
        N576, N575, N574, N573}) );
  FPU_CAL_DW01_inc_3 add_175 ( .A({n285, E[7:0]}), .SUM({N513, N512, N511, 
        N510, N509, N508, N507, N506, N505}) );
  FPU_CAL_DW01_add_0 add_117 ( .A({1'b0, n65, A[29:23]}), .B({1'b0, N437, 
        B[29:24], n31}), .CI(1'b0), .SUM({N338, N337, N336, N335, N334, N333, 
        N332, N331, N330}) );
  FPU_CAL_DW01_sub_2 sub_88 ( .A({1'b0, N134, N133, N132, N131, N130, N129, 
        N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, 
        N116, N115, N114, N113, N112, N111}), .B({1'b0, N166, N165, N164, N163, 
        N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, 
        N150, N149, N148, N147, N146, N145, N144, N143}), .CI(1'b0), .DIFF({
        N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, 
        N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, 
        N248}) );
  FPU_CAL_DW01_sub_3 sub_82 ( .A({1'b0, N166, N165, N164, N163, N162, N161, 
        N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, 
        N148, N147, N146, N145, N144, N143}), .B({1'b0, N134, N133, N132, N131, 
        N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, 
        N118, N117, N116, N115, N114, N113, N112, N111}), .CI(1'b0), .DIFF({
        N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, 
        N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, 
        N172}) );
  FPU_CAL_DW01_add_1 r226 ( .A({1'b0, N166, N165, N164, N163, N162, N161, N160, 
        N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, 
        N147, N146, N145, N144, N143}), .B({1'b0, N134, N133, N132, N131, N130, 
        N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, 
        N117, N116, N115, N114, N113, N112, N111}), .CI(1'b0), .SUM({N221, 
        N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, 
        N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197}) );
  FPU_CAL_DW_rash_0 srl_75 ( .A({1'b1, n139, A[21], n136, n132, A[18:16], n122, 
        A[14:0]}), .DATA_TC(1'b0), .SH({N86, N85, N84, N83, N82, N81, N80, N79}), .SH_TC(1'b0), .B({N110, N109, N108, N107, N106, N105, N104, N103, N102, 
        N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, 
        N87}) );
  FPU_CAL_DW01_sub_4 sub_75 ( .A({N437, B[29:24], n32}), .B({n65, A[29:23]}), 
        .CI(1'b0), .DIFF({N86, N85, N84, N83, N82, N81, N80, N79}) );
  FPU_CAL_DW_rash_1 srl_71 ( .A({1'b1, B[22:0]}), .DATA_TC(1'b0), .SH({N54, 
        N53, N52, N51, N50, N49, N48, N47}), .SH_TC(1'b0), .B({N78, N77, N76, 
        N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, 
        N61, N60, N59, N58, N57, N56, N55}) );
  FPU_CAL_DW01_sub_5 sub_71 ( .A({n65, A[29:23]}), .B({N437, B[29:24], n31}), 
        .CI(1'b0), .DIFF({N54, N53, N52, N51, N50, N49, N48, N47}) );
  FPU_CAL_DW01_add_4 add_0_root_sub_0_root_sub_122 ( .A({1'b0, n65, A[29:23]}), 
        .B({n43, N350, N349, N348, N347, N346, N345, N344, n55}), .CI(1'b0), 
        .SUM({N360, N359, N358, N357, N356, N355, N354, N353, N352}) );
  FPU_CAL_DW02_mult_0 mult_123 ( .A({1'b1, n139, A[21], n136, n132, A[18:16], 
        n122, A[14:0]}), .B({1'b1, B[22:0]}), .TC(1'b0), .PRODUCT({N408, N407, 
        N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, 
        N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, 
        N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, 
        N370, N369, N368, N367, N366, N365, N364, N363, N362, N361}) );
  FPU_CAL_DW01_add_3 add_0_root_sub_0_root_add_150 ( .A({1'b0, n65, A[29:23]}), 
        .B({N437, N437, n59, n654, n58, n57, n56, n653, n55}), .CI(1'b0), 
        .SUM({N446, N445, N444, N443, N442, N441, N440, N439, N438}) );
  FPU_CAL_DW01_inc_4 add_0_root_add_170 ( .A({N492, N491, N490, N489, N488, 
        N487, N486, N485, N484}), .SUM({N501, N500, N499, N498, N497, N496, 
        N495, N494, N493}) );
  FPU_CAL_DW_div_uns_2 r243 ( .a({1'b1, div[46:25], n22, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({1'b1, 
        divider[22:2], n24, divider[0]}), .quotient({SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, N536, N527, N526, N525, N524, N523, N522, 
        N521, N520, N519, SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, 
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52}) );
  DFFX1_RVT \M_sum_reg[8]  ( .D(n45), .CLK(clk), .Q(M_sum[8]), .QN(n729) );
  DFFX1_RVT \M1M2_reg[40]  ( .D(n432), .CLK(clk), .Q(M1M2[40]) );
  DFFX1_RVT \M1M2_reg[41]  ( .D(n431), .CLK(clk), .Q(M1M2[41]) );
  DFFX1_RVT \M1M2_reg[42]  ( .D(n430), .CLK(clk), .Q(M1M2[42]) );
  DFFX1_RVT \M1M2_reg[43]  ( .D(n429), .CLK(clk), .Q(M1M2[43]) );
  DFFX1_RVT \M1M2_reg[44]  ( .D(n428), .CLK(clk), .Q(M1M2[44]) );
  DFFX1_RVT \M1M2_reg[45]  ( .D(n427), .CLK(clk), .Q(M1M2[45]) );
  DFFX1_RVT \M1M2_reg[39]  ( .D(n433), .CLK(clk), .Q(M1M2[39]) );
  DFFX1_RVT \quotient_reg[18]  ( .D(n395), .CLK(clk), .Q(quotient[18]) );
  DFFX1_RVT \quotient_reg[17]  ( .D(n394), .CLK(clk), .Q(quotient[17]) );
  DFFX1_RVT \M1M2_reg[46]  ( .D(n426), .CLK(clk), .Q(M1M2[46]) );
  DFFX1_RVT \quotient_reg[15]  ( .D(n392), .CLK(clk), .Q(quotient[15]) );
  DFFX1_RVT \quotient_reg[16]  ( .D(n393), .CLK(clk), .Q(quotient[16]) );
  DFFX1_RVT \E_reg[6]  ( .D(n524), .CLK(clk), .Q(E[6]), .QN(n742) );
  DFFX1_RVT \E_reg[0]  ( .D(n530), .CLK(clk), .Q(E[0]), .QN(n738) );
  DFFX1_RVT \E_reg[5]  ( .D(n525), .CLK(clk), .Q(E[5]), .QN(n140) );
  DFFX1_RVT \E_reg[7]  ( .D(n523), .CLK(clk), .Q(E[7]), .QN(n740) );
  DFFX1_RVT \E_reg[4]  ( .D(n526), .CLK(clk), .Q(E[4]), .QN(n141) );
  DFFX1_RVT \E_reg[2]  ( .D(n528), .CLK(clk), .Q(E[2]), .QN(n743) );
  DFFX1_RVT \E_reg[3]  ( .D(n527), .CLK(clk), .Q(E[3]), .QN(n744) );
  DFFX1_RVT \E_reg[1]  ( .D(n529), .CLK(clk), .Q(E[1]), .QN(n739) );
  DFFX1_RVT \M_sum_reg[4]  ( .D(n517), .CLK(clk), .Q(n260), .QN(n727) );
  DFFX1_RVT \M_sum_reg[2]  ( .D(n18), .CLK(clk), .Q(n264), .QN(n714) );
  DFFX1_RVT \M_sum_reg[3]  ( .D(n518), .CLK(clk), .Q(n262), .QN(n725) );
  DFFX1_RVT \M_sum_reg[1]  ( .D(n520), .CLK(clk), .Q(n266), .QN(n719) );
  DFFX1_RVT \M_sum_reg[18]  ( .D(n503), .CLK(clk), .Q(n241), .QN(n718) );
  DFFX1_RVT \M_sum_reg[22]  ( .D(n14), .CLK(clk), .Q(n233), .QN(n723) );
  DFFX1_RVT \M_sum_reg[19]  ( .D(n13), .CLK(clk), .Q(n239), .QN(n720) );
  DFFX1_RVT \M_sum_reg[23]  ( .D(n498), .CLK(clk), .Q(n231), .QN(n713) );
  DFFX1_RVT \M_sum_reg[24]  ( .D(n497), .CLK(clk), .Q(n229), .QN(n715) );
  DFFX1_RVT \M_sum_reg[20]  ( .D(n501), .CLK(clk), .Q(n237), .QN(n722) );
  DFFX1_RVT \M_sum_reg[17]  ( .D(n504), .CLK(clk), .Q(n243), .QN(n736) );
  DFFX1_RVT \M_sum_reg[21]  ( .D(n500), .CLK(clk), .Q(n235), .QN(n724) );
  DFFX1_RVT \M_sum_reg[9]  ( .D(n512), .CLK(clk), .Q(n254), .QN(n728) );
  DFFX1_RVT \M_sum_reg[16]  ( .D(n505), .CLK(clk), .Q(n245), .QN(n737) );
  DFFX1_RVT \divider_reg[1]  ( .D(n494), .CLK(clk), .Q(divider[1]), .QN(n23)
         );
  DFFX1_RVT \M_sum_reg[0]  ( .D(n17), .CLK(clk), .Q(n268), .QN(n732) );
  DFFX1_RVT \M1M2_reg[0]  ( .D(n472), .CLK(clk), .Q(n184) );
  DFFX1_RVT \M1M2_reg[8]  ( .D(n464), .CLK(clk), .Q(n192) );
  DFFX1_RVT \M1M2_reg[7]  ( .D(n465), .CLK(clk), .Q(n191) );
  DFFX1_RVT \M1M2_reg[6]  ( .D(n466), .CLK(clk), .Q(n190) );
  DFFX1_RVT \M1M2_reg[5]  ( .D(n467), .CLK(clk), .Q(n189) );
  DFFX1_RVT \M1M2_reg[4]  ( .D(n468), .CLK(clk), .Q(n188) );
  DFFX1_RVT \M1M2_reg[3]  ( .D(n469), .CLK(clk), .Q(n187) );
  DFFX1_RVT \M1M2_reg[2]  ( .D(n470), .CLK(clk), .Q(n186) );
  DFFX1_RVT \M1M2_reg[1]  ( .D(n471), .CLK(clk), .Q(n185) );
  DFFX1_RVT \M1M2_reg[9]  ( .D(n463), .CLK(clk), .Q(n193) );
  DFFX1_RVT \M1M2_reg[10]  ( .D(n462), .CLK(clk), .Q(n194) );
  DFFX1_RVT \M1M2_reg[11]  ( .D(n461), .CLK(clk), .Q(n195) );
  DFFX1_RVT \M1M2_reg[12]  ( .D(n460), .CLK(clk), .Q(n196) );
  DFFX1_RVT \M1M2_reg[13]  ( .D(n459), .CLK(clk), .Q(n197) );
  DFFX1_RVT \M1M2_reg[14]  ( .D(n458), .CLK(clk), .Q(n198) );
  DFFX1_RVT \M1M2_reg[15]  ( .D(n457), .CLK(clk), .Q(n199) );
  DFFX1_RVT \M1M2_reg[16]  ( .D(n456), .CLK(clk), .Q(n200) );
  DFFX1_RVT \M1M2_reg[17]  ( .D(n455), .CLK(clk), .Q(n201) );
  DFFX1_RVT \M1M2_reg[18]  ( .D(n454), .CLK(clk), .Q(n203) );
  DFFX1_RVT \M1M2_reg[19]  ( .D(n453), .CLK(clk), .Q(n204) );
  DFFX1_RVT \M1M2_reg[20]  ( .D(n452), .CLK(clk), .Q(n205) );
  DFFX1_RVT \M1M2_reg[21]  ( .D(n451), .CLK(clk), .Q(n206) );
  DFFX1_RVT \M1M2_reg[22]  ( .D(n450), .CLK(clk), .Q(n207) );
  DFFX1_RVT \M1M2_reg[23]  ( .D(n449), .CLK(clk), .Q(n208) );
  DFFX1_RVT \M1M2_reg[24]  ( .D(n448), .CLK(clk), .Q(n209) );
  DFFX1_RVT \M1M2_reg[25]  ( .D(n447), .CLK(clk), .Q(n210) );
  DFFX1_RVT \M1M2_reg[26]  ( .D(n446), .CLK(clk), .Q(n212) );
  DFFX1_RVT \M1M2_reg[27]  ( .D(n445), .CLK(clk), .Q(n213) );
  DFFX1_RVT \M1M2_reg[28]  ( .D(n444), .CLK(clk), .Q(n215) );
  DFFX1_RVT \M1M2_reg[29]  ( .D(n443), .CLK(clk), .Q(n216) );
  DFFX1_RVT \M1M2_reg[30]  ( .D(n442), .CLK(clk), .Q(n218) );
  DFFX1_RVT \M1M2_reg[31]  ( .D(n441), .CLK(clk), .Q(n219) );
  DFFX1_RVT \M1M2_reg[32]  ( .D(n440), .CLK(clk), .Q(n221) );
  DFFX1_RVT \M1M2_reg[33]  ( .D(n439), .CLK(clk), .Q(n222) );
  DFFX1_RVT \M1M2_reg[34]  ( .D(n438), .CLK(clk), .Q(n224) );
  DFFX1_RVT \M1M2_reg[35]  ( .D(n437), .CLK(clk), .Q(n225) );
  DFFX1_RVT \M1M2_reg[36]  ( .D(n436), .CLK(clk), .Q(n227) );
  DFFX1_RVT \M1M2_reg[37]  ( .D(n435), .CLK(clk), .Q(n228) );
  DFFX1_RVT \M1M2_reg[38]  ( .D(n434), .CLK(clk), .Q(n287) );
  DFFX1_RVT \M1M2_reg[47]  ( .D(n531), .CLK(clk), .Q(n279), .QN(n143) );
  DFFX1_RVT error_reg ( .D(n425), .CLK(clk), .Q(error) );
  DFFX1_RVT \div_reg[38]  ( .D(n415), .CLK(clk), .Q(div[38]) );
  DFFX1_RVT \div_reg[43]  ( .D(n420), .CLK(clk), .Q(div[43]) );
  DFFX1_RVT \div_reg[46]  ( .D(n423), .CLK(clk), .Q(div[46]) );
  DFFX1_RVT \div_reg[41]  ( .D(n418), .CLK(clk), .Q(div[41]) );
  DFFX1_RVT \div_reg[39]  ( .D(n416), .CLK(clk), .Q(div[39]) );
  DFFX1_RVT \div_reg[42]  ( .D(n419), .CLK(clk), .Q(div[42]) );
  DFFX1_RVT \div_reg[37]  ( .D(n414), .CLK(clk), .Q(div[37]) );
  DFFX1_RVT \div_reg[40]  ( .D(n417), .CLK(clk), .Q(div[40]) );
  DFFX1_RVT \div_reg[45]  ( .D(n422), .CLK(clk), .Q(div[45]) );
  DFFX1_RVT \div_reg[44]  ( .D(n421), .CLK(clk), .Q(div[44]) );
  DFFX1_RVT over_flow_reg ( .D(n424), .CLK(clk), .Q(over_flow) );
  DFFX1_RVT \next_state_reg[1]  ( .D(n522), .CLK(clk), .Q(next_state[1]), .QN(
        n291) );
  DFFX1_RVT \divider_reg[22]  ( .D(n473), .CLK(clk), .Q(divider[22]) );
  DFFX1_RVT \divider_reg[21]  ( .D(n474), .CLK(clk), .Q(divider[21]) );
  DFFX1_RVT \divider_reg[20]  ( .D(n475), .CLK(clk), .Q(divider[20]) );
  DFFX1_RVT \divider_reg[19]  ( .D(n476), .CLK(clk), .Q(divider[19]) );
  DFFX1_RVT \divider_reg[18]  ( .D(n477), .CLK(clk), .Q(divider[18]) );
  DFFX1_RVT \divider_reg[17]  ( .D(n478), .CLK(clk), .Q(divider[17]) );
  DFFX1_RVT \divider_reg[16]  ( .D(n479), .CLK(clk), .Q(divider[16]) );
  DFFX1_RVT \divider_reg[15]  ( .D(n480), .CLK(clk), .Q(divider[15]) );
  DFFX1_RVT \divider_reg[14]  ( .D(n481), .CLK(clk), .Q(divider[14]) );
  DFFX1_RVT \divider_reg[13]  ( .D(n482), .CLK(clk), .Q(divider[13]) );
  DFFX1_RVT \divider_reg[12]  ( .D(n483), .CLK(clk), .Q(divider[12]) );
  DFFX1_RVT \divider_reg[11]  ( .D(n484), .CLK(clk), .Q(divider[11]) );
  DFFX1_RVT \divider_reg[10]  ( .D(n485), .CLK(clk), .Q(divider[10]) );
  DFFX1_RVT \divider_reg[9]  ( .D(n486), .CLK(clk), .Q(divider[9]) );
  DFFX1_RVT \divider_reg[8]  ( .D(n487), .CLK(clk), .Q(divider[8]) );
  DFFX1_RVT \divider_reg[7]  ( .D(n488), .CLK(clk), .Q(divider[7]) );
  DFFX1_RVT \divider_reg[6]  ( .D(n489), .CLK(clk), .Q(divider[6]) );
  DFFX1_RVT \divider_reg[5]  ( .D(n490), .CLK(clk), .Q(divider[5]) );
  DFFX1_RVT \divider_reg[4]  ( .D(n491), .CLK(clk), .Q(divider[4]) );
  DFFX1_RVT \divider_reg[3]  ( .D(n492), .CLK(clk), .Q(divider[3]) );
  DFFX1_RVT \divider_reg[2]  ( .D(n493), .CLK(clk), .Q(divider[2]) );
  DFFX1_RVT \divider_reg[0]  ( .D(n495), .CLK(clk), .Q(divider[0]) );
  DFFX1_RVT \div_reg[36]  ( .D(n413), .CLK(clk), .Q(div[36]) );
  DFFX1_RVT \div_reg[35]  ( .D(n412), .CLK(clk), .Q(div[35]) );
  DFFX1_RVT \div_reg[34]  ( .D(n411), .CLK(clk), .Q(div[34]) );
  DFFX1_RVT \div_reg[33]  ( .D(n410), .CLK(clk), .Q(div[33]) );
  DFFX1_RVT \div_reg[32]  ( .D(n409), .CLK(clk), .Q(div[32]) );
  DFFX1_RVT \div_reg[31]  ( .D(n408), .CLK(clk), .Q(div[31]) );
  DFFX1_RVT \div_reg[30]  ( .D(n407), .CLK(clk), .Q(div[30]) );
  DFFX1_RVT \div_reg[29]  ( .D(n406), .CLK(clk), .Q(div[29]) );
  DFFX1_RVT \div_reg[28]  ( .D(n405), .CLK(clk), .Q(div[28]) );
  DFFX1_RVT \div_reg[27]  ( .D(n404), .CLK(clk), .Q(div[27]) );
  DFFX1_RVT \div_reg[26]  ( .D(n403), .CLK(clk), .Q(div[26]) );
  DFFX1_RVT \div_reg[25]  ( .D(n402), .CLK(clk), .Q(div[25]) );
  DFFX1_RVT \next_state_reg[0]  ( .D(n532), .CLK(clk), .Q(next_state[0]), .QN(
        n581) );
  DFFX1_RVT \Y_reg[31]  ( .D(n382), .CLK(clk), .Q(Y[31]) );
  DFFX1_RVT \Y_reg[30]  ( .D(n383), .CLK(clk), .Q(Y[30]) );
  DFFX1_RVT \Y_reg[29]  ( .D(n384), .CLK(clk), .Q(Y[29]) );
  DFFX1_RVT \Y_reg[28]  ( .D(n385), .CLK(clk), .Q(Y[28]) );
  DFFX1_RVT \Y_reg[27]  ( .D(n386), .CLK(clk), .Q(Y[27]) );
  DFFX1_RVT \Y_reg[26]  ( .D(n387), .CLK(clk), .Q(Y[26]) );
  DFFX1_RVT \Y_reg[25]  ( .D(n388), .CLK(clk), .Q(Y[25]) );
  DFFX1_RVT \Y_reg[24]  ( .D(n389), .CLK(clk), .Q(Y[24]) );
  DFFX1_RVT \Y_reg[23]  ( .D(n390), .CLK(clk), .Q(Y[23]) );
  DFFX1_RVT \Y_reg[22]  ( .D(n391), .CLK(clk), .Q(Y[22]) );
  DFFX1_RVT \quotient_reg[23]  ( .D(n400), .CLK(clk), .Q(quotient[23]) );
  DFFX1_RVT S_reg ( .D(n496), .CLK(clk), .Q(n564) );
  DFFX1_RVT \quotient_reg[22]  ( .D(n399), .CLK(clk), .Q(quotient[22]) );
  DFFX1_RVT \quotient_reg[21]  ( .D(n398), .CLK(clk), .Q(quotient[21]) );
  DFFX1_RVT \quotient_reg[20]  ( .D(n397), .CLK(clk), .Q(quotient[20]) );
  DFFX1_RVT \quotient_reg[19]  ( .D(n396), .CLK(clk), .Q(quotient[19]) );
  DFFX1_RVT \M_sum_reg[15]  ( .D(n506), .CLK(clk), .Q(M_sum[15]), .QN(n735) );
  DFFX1_RVT \M_sum_reg[14]  ( .D(n507), .CLK(clk), .Q(n288), .QN(n721) );
  DFFX1_RVT \M_sum_reg[13]  ( .D(n15), .CLK(clk), .Q(n247), .QN(n717) );
  DFFX1_RVT \M_sum_reg[12]  ( .D(n509), .CLK(clk), .Q(n249), .QN(n716) );
  DFFX1_RVT \M_sum_reg[11]  ( .D(n510), .CLK(clk), .Q(n251), .QN(n733) );
  DFFX1_RVT \M_sum_reg[10]  ( .D(n511), .CLK(clk), .Q(n252), .QN(n734) );
  DFFX1_RVT \M_sum_reg[6]  ( .D(n515), .CLK(clk), .Q(n256), .QN(n731) );
  DFFX1_RVT \M_sum_reg[5]  ( .D(n516), .CLK(clk), .Q(n258), .QN(n726) );
  DFFX1_RVT \M_sum_reg[7]  ( .D(n514), .CLK(clk), .Q(n255), .QN(n730) );
  DFFX1_RVT \div_reg[24]  ( .D(n401), .CLK(clk), .Q(div[24]), .QN(n21) );
  INVX1_RVT U3 ( .A(n21), .Y(n22) );
  INVX1_RVT U5 ( .A(N122), .Y(n340) );
  INVX1_RVT U7 ( .A(N123), .Y(n339) );
  INVX1_RVT U9 ( .A(N125), .Y(n332) );
  INVX1_RVT U11 ( .A(N126), .Y(n337) );
  OA21X1_RVT U13 ( .A1(A[24]), .A2(n653), .A3(n55), .Y(n712) );
  AND4X1_RVT U15 ( .A1(A[27]), .A2(A[26]), .A3(A[25]), .A4(A[24]), .Y(n679) );
  INVX1_RVT U58 ( .A(A[24]), .Y(n650) );
  INVX1_RVT U60 ( .A(N133), .Y(n325) );
  INVX1_RVT U61 ( .A(n619), .Y(n626) );
  INVX1_RVT U62 ( .A(A[20]), .Y(n137) );
  INVX1_RVT U63 ( .A(A[22]), .Y(n142) );
  INVX1_RVT U64 ( .A(A[19]), .Y(n134) );
  MUX21X1_RVT U65 ( .A1(N90), .A2(A[3]), .S0(n88), .Y(N146) );
  INVX1_RVT U66 ( .A(n281), .Y(n180) );
  MUX21X1_RVT U67 ( .A1(N95), .A2(A[8]), .S0(n89), .Y(N151) );
  NAND2X0_RVT U68 ( .A1(N259), .A2(n86), .Y(n29) );
  INVX1_RVT U69 ( .A(N185), .Y(n26) );
  INVX1_RVT U70 ( .A(N261), .Y(n25) );
  INVX1_RVT U71 ( .A(n50), .Y(n512) );
  AO221X1_RVT U72 ( .A1(N196), .A2(n82), .A3(N272), .A4(n85), .A5(n230), .Y(
        n497) );
  NAND2X0_RVT U73 ( .A1(n6), .A2(n19), .Y(n510) );
  NOR2X1_RVT U74 ( .A1(n9), .A2(n26), .Y(n28) );
  INVX1_RVT U75 ( .A(A[8]), .Y(n114) );
  NAND3X0_RVT U76 ( .A1(n40), .A2(n176), .A3(n563), .Y(n1) );
  INVX1_RVT U77 ( .A(A[9]), .Y(n115) );
  AND3X1_RVT U78 ( .A1(n558), .A2(n376), .A3(n11), .Y(n2) );
  INVX1_RVT U79 ( .A(A[10]), .Y(n116) );
  AND2X1_RVT U80 ( .A1(N134), .A2(n8), .Y(n3) );
  OAI22X1_RVT U81 ( .A1(n16), .A2(n44), .A3(n40), .A4(n729), .Y(n4) );
  OAI22X1_RVT U82 ( .A1(n33), .A2(n16), .A3(n40), .A4(n728), .Y(n5) );
  MUX21X1_RVT U83 ( .A1(N99), .A2(A[12]), .S0(n91), .Y(N155) );
  MUX21X1_RVT U84 ( .A1(A[0]), .A2(N87), .S0(n101), .Y(N143) );
  AOI22X1_RVT U85 ( .A1(N208), .A2(n83), .A3(n103), .A4(n251), .Y(n6) );
  OAI22X1_RVT U86 ( .A1(n51), .A2(n16), .A3(n40), .A4(n735), .Y(n7) );
  AOI21X1_RVT U87 ( .A1(N165), .A2(n325), .A3(n318), .Y(n8) );
  NAND3X0_RVT U88 ( .A1(n563), .A2(N167), .A3(n40), .Y(n9) );
  AND2X1_RVT U89 ( .A1(n297), .A2(n289), .Y(n10) );
  AND2X1_RVT U90 ( .A1(n147), .A2(n291), .Y(n11) );
  INVX1_RVT U91 ( .A(A[6]), .Y(n112) );
  INVX1_RVT U92 ( .A(A[21]), .Y(n138) );
  OR2X1_RVT U93 ( .A1(n27), .A2(n28), .Y(n12) );
  AO221X1_RVT U94 ( .A1(N191), .A2(n82), .A3(N267), .A4(n85), .A5(n240), .Y(
        n13) );
  AO221X1_RVT U95 ( .A1(N194), .A2(n82), .A3(N270), .A4(n85), .A5(n234), .Y(
        n14) );
  OR2X1_RVT U96 ( .A1(n248), .A2(n12), .Y(n15) );
  MUX21X1_RVT U97 ( .A1(N94), .A2(A[7]), .S0(n89), .Y(N150) );
  NAND2X0_RVT U98 ( .A1(n567), .A2(n40), .Y(n16) );
  OAI221X1_RVT U99 ( .A1(n34), .A2(n9), .A3(n35), .A4(n48), .A5(n36), .Y(n17)
         );
  AO221X1_RVT U100 ( .A1(N184), .A2(n82), .A3(N260), .A4(n86), .A5(n250), .Y(
        n509) );
  AO221X1_RVT U101 ( .A1(N174), .A2(n81), .A3(N250), .A4(n86), .A5(n265), .Y(
        n18) );
  AND2X1_RVT U102 ( .A1(n29), .A2(n30), .Y(n19) );
  AND4X1_RVT U103 ( .A1(n696), .A2(n375), .A3(n290), .A4(n282), .Y(n20) );
  INVX1_RVT U104 ( .A(n280), .Y(n179) );
  INVX1_RVT U105 ( .A(n23), .Y(n24) );
  MUX21X1_RVT U106 ( .A1(N102), .A2(n122), .S0(n93), .Y(N158) );
  NOR2X1_RVT U107 ( .A1(n48), .A2(n25), .Y(n27) );
  NAND2X0_RVT U108 ( .A1(N183), .A2(n81), .Y(n30) );
  INVX1_RVT U109 ( .A(n1), .Y(n85) );
  INVX1_RVT U110 ( .A(n560), .Y(n96) );
  INVX1_RVT U111 ( .A(n86), .Y(n48) );
  INVX1_RVT U112 ( .A(n55), .Y(n32) );
  INVX1_RVT U113 ( .A(n55), .Y(n31) );
  INVX1_RVT U114 ( .A(N172), .Y(n34) );
  INVX1_RVT U115 ( .A(N248), .Y(n35) );
  INVX1_RVT U116 ( .A(n64), .Y(n65) );
  INVX1_RVT U117 ( .A(A[30]), .Y(n64) );
  INVX1_RVT U118 ( .A(A[5]), .Y(n111) );
  INVX1_RVT U119 ( .A(A[7]), .Y(n113) );
  INVX1_RVT U120 ( .A(A[13]), .Y(n119) );
  INVX1_RVT U121 ( .A(A[15]), .Y(n124) );
  INVX1_RVT U122 ( .A(A[17]), .Y(n128) );
  INVX1_RVT U123 ( .A(A[16]), .Y(n126) );
  INVX1_RVT U124 ( .A(A[12]), .Y(n118) );
  INVX1_RVT U125 ( .A(A[4]), .Y(n110) );
  INVX1_RVT U126 ( .A(A[14]), .Y(n120) );
  INVX1_RVT U127 ( .A(A[18]), .Y(n130) );
  INVX1_RVT U128 ( .A(N206), .Y(n33) );
  INVX0_RVT U129 ( .A(n40), .Y(n103) );
  INVX0_RVT U130 ( .A(N120), .Y(n330) );
  INVX0_RVT U131 ( .A(N119), .Y(n331) );
  INVX0_RVT U132 ( .A(N116), .Y(n335) );
  INVX0_RVT U133 ( .A(N114), .Y(n319) );
  INVX1_RVT U134 ( .A(N166), .Y(n38) );
  INVX1_RVT U135 ( .A(A[28]), .Y(n62) );
  INVX1_RVT U136 ( .A(B[29]), .Y(n59) );
  INVX0_RVT U137 ( .A(n9), .Y(n82) );
  NOR4X1_RVT U138 ( .A1(n607), .A2(n631), .A3(n622), .A4(n621), .Y(n634) );
  AOI22X1_RVT U139 ( .A1(N197), .A2(n83), .A3(n103), .A4(n268), .Y(n36) );
  INVX1_RVT U140 ( .A(N121), .Y(n341) );
  INVX1_RVT U141 ( .A(N115), .Y(n336) );
  INVX1_RVT U142 ( .A(N124), .Y(n338) );
  INVX1_RVT U143 ( .A(N118), .Y(n333) );
  INVX1_RVT U144 ( .A(N132), .Y(n322) );
  OAI221X1_RVT U145 ( .A1(n52), .A2(N131), .A3(n53), .A4(N132), .A5(n54), .Y(
        n37) );
  INVX1_RVT U146 ( .A(A[25]), .Y(n60) );
  INVX1_RVT U147 ( .A(A[29]), .Y(n63) );
  INVX1_RVT U148 ( .A(B[25]), .Y(n56) );
  INVX1_RVT U149 ( .A(n280), .Y(n66) );
  INVX1_RVT U150 ( .A(n280), .Y(n67) );
  INVX1_RVT U151 ( .A(n280), .Y(n68) );
  INVX1_RVT U152 ( .A(n94), .Y(n101) );
  INVX1_RVT U153 ( .A(n95), .Y(n102) );
  INVX1_RVT U154 ( .A(n96), .Y(n94) );
  INVX1_RVT U155 ( .A(n98), .Y(n91) );
  INVX1_RVT U156 ( .A(n98), .Y(n92) );
  INVX1_RVT U157 ( .A(n97), .Y(n93) );
  INVX1_RVT U158 ( .A(N164), .Y(n53) );
  INVX1_RVT U159 ( .A(n96), .Y(n95) );
  INVX1_RVT U160 ( .A(n99), .Y(n89) );
  INVX1_RVT U161 ( .A(n99), .Y(n88) );
  INVX1_RVT U162 ( .A(n98), .Y(n90) );
  INVX1_RVT U163 ( .A(n16), .Y(n83) );
  INVX1_RVT U164 ( .A(n16), .Y(n84) );
  INVX1_RVT U165 ( .A(shifted[0]), .Y(n105) );
  INVX1_RVT U166 ( .A(n574), .Y(n289) );
  OAI22X1_RVT U167 ( .A1(n8), .A2(N134), .A3(n38), .A4(n3), .Y(N167) );
  INVX0_RVT U168 ( .A(N212), .Y(n51) );
  INVX0_RVT U169 ( .A(n560), .Y(n98) );
  INVX1_RVT U170 ( .A(n560), .Y(n97) );
  INVX0_RVT U171 ( .A(n560), .Y(n99) );
  INVX1_RVT U172 ( .A(n100), .Y(n87) );
  INVX1_RVT U173 ( .A(n560), .Y(n100) );
  INVX1_RVT U174 ( .A(\sub_1_root_add_170/carry[7] ), .Y(n283) );
  INVX1_RVT U175 ( .A(n576), .Y(n369) );
  AND2X1_RVT U176 ( .A1(n559), .A2(n290), .Y(n519) );
  AND2X1_RVT U177 ( .A1(n568), .A2(n558), .Y(n513) );
  AND2X1_RVT U178 ( .A1(n559), .A2(n561), .Y(n368) );
  INVX1_RVT U179 ( .A(n277), .Y(n174) );
  INVX1_RVT U180 ( .A(n171), .Y(n170) );
  INVX1_RVT U181 ( .A(n40), .Y(n104) );
  NAND2X0_RVT U182 ( .A1(n11), .A2(n290), .Y(n574) );
  INVX1_RVT U183 ( .A(n183), .Y(n71) );
  INVX1_RVT U184 ( .A(n183), .Y(n70) );
  INVX1_RVT U185 ( .A(n183), .Y(n69) );
  INVX1_RVT U186 ( .A(n183), .Y(n72) );
  INVX1_RVT U187 ( .A(n181), .Y(n79) );
  INVX1_RVT U188 ( .A(n181), .Y(n78) );
  INVX1_RVT U189 ( .A(n181), .Y(n77) );
  INVX1_RVT U190 ( .A(n181), .Y(n80) );
  INVX1_RVT U191 ( .A(n182), .Y(n73) );
  INVX1_RVT U192 ( .A(n182), .Y(n74) );
  INVX1_RVT U193 ( .A(n182), .Y(n75) );
  INVX1_RVT U194 ( .A(n182), .Y(n76) );
  AND3X1_RVT U195 ( .A1(n594), .A2(n375), .A3(n290), .Y(n39) );
  INVX1_RVT U196 ( .A(N205), .Y(n44) );
  AND3X1_RVT U197 ( .A1(n660), .A2(n376), .A3(n292), .Y(n40) );
  INVX1_RVT U198 ( .A(n134), .Y(n132) );
  INVX1_RVT U199 ( .A(n124), .Y(n122) );
  INVX1_RVT U200 ( .A(n137), .Y(n136) );
  INVX1_RVT U201 ( .A(n608), .Y(n290) );
  INVX1_RVT U202 ( .A(N163), .Y(n52) );
  AO221X1_RVT U203 ( .A1(N151), .A2(n331), .A3(N152), .A4(n330), .A5(n306), 
        .Y(n307) );
  AO221X1_RVT U204 ( .A1(N159), .A2(n329), .A3(N160), .A4(n328), .A5(n314), 
        .Y(n315) );
  INVX1_RVT U205 ( .A(N127), .Y(n329) );
  INVX1_RVT U206 ( .A(N130), .Y(n326) );
  INVX1_RVT U207 ( .A(N255), .Y(n47) );
  INVX1_RVT U208 ( .A(N128), .Y(n328) );
  INVX1_RVT U209 ( .A(N112), .Y(n321) );
  INVX1_RVT U210 ( .A(N131), .Y(n324) );
  INVX1_RVT U211 ( .A(N129), .Y(n327) );
  INVX1_RVT U212 ( .A(N113), .Y(n320) );
  INVX1_RVT U213 ( .A(N117), .Y(n334) );
  INVX0_RVT U214 ( .A(n284), .Y(n146) );
  AND2X1_RVT U215 ( .A1(n577), .A2(n576), .Y(n596) );
  INVX1_RVT U216 ( .A(n159), .Y(n158) );
  AND2X1_RVT U217 ( .A1(N516), .A2(n289), .Y(n41) );
  INVX1_RVT U218 ( .A(n151), .Y(n150) );
  INVX1_RVT U219 ( .A(n167), .Y(n166) );
  INVX1_RVT U220 ( .A(N516), .Y(n297) );
  INVX1_RVT U221 ( .A(n607), .Y(n561) );
  OR3X2_RVT U222 ( .A1(n367), .A2(N338), .A3(N337), .Y(n42) );
  INVX1_RVT U223 ( .A(n380), .Y(n147) );
  INVX1_RVT U224 ( .A(n697), .Y(n282) );
  INVX1_RVT U225 ( .A(n163), .Y(n162) );
  NOR2X0_RVT U226 ( .A1(N437), .A2(\sub_1_root_sub_0_root_sub_122/carry[7] ), 
        .Y(n43) );
  INVX1_RVT U227 ( .A(start), .Y(n144) );
  INVX1_RVT U228 ( .A(A[26]), .Y(n61) );
  INVX1_RVT U229 ( .A(B[27]), .Y(n58) );
  INVX1_RVT U230 ( .A(B[26]), .Y(n57) );
  INVX1_RVT U231 ( .A(A[1]), .Y(n107) );
  INVX1_RVT U232 ( .A(A[3]), .Y(n109) );
  INVX1_RVT U233 ( .A(A[2]), .Y(n108) );
  INVX1_RVT U234 ( .A(A[0]), .Y(n106) );
  AO221X1_RVT U235 ( .A1(N173), .A2(n81), .A3(N249), .A4(n86), .A5(n267), .Y(
        n520) );
  FADDX1_RVT U236 ( .A(E[1]), .B(n296), .CI(\sub_1_root_add_170/carry[1] ), 
        .CO(\sub_1_root_add_170/carry[2] ), .S(N485) );
  INVX1_RVT U237 ( .A(shifted[1]), .Y(n296) );
  FADDX1_RVT U238 ( .A(E[4]), .B(n293), .CI(\sub_1_root_add_170/carry[4] ), 
        .CO(\sub_1_root_add_170/carry[5] ), .S(N488) );
  INVX1_RVT U239 ( .A(shifted[4]), .Y(n293) );
  FADDX1_RVT U240 ( .A(E[2]), .B(n295), .CI(\sub_1_root_add_170/carry[2] ), 
        .CO(\sub_1_root_add_170/carry[3] ), .S(N486) );
  INVX1_RVT U241 ( .A(shifted[2]), .Y(n295) );
  FADDX1_RVT U242 ( .A(E[3]), .B(n294), .CI(\sub_1_root_add_170/carry[3] ), 
        .CO(\sub_1_root_add_170/carry[4] ), .S(N487) );
  INVX1_RVT U243 ( .A(shifted[3]), .Y(n294) );
  XNOR2X1_RVT U244 ( .A1(n278), .A2(n285), .Y(N545) );
  AO21X1_RVT U245 ( .A1(E[6]), .A2(n171), .A3(n174), .Y(n173) );
  OR2X1_RVT U246 ( .A1(E[7]), .A2(n277), .Y(n278) );
  INVX1_RVT U247 ( .A(A[23]), .Y(n648) );
  INVX1_RVT U248 ( .A(B[23]), .Y(n55) );
  INVX1_RVT U249 ( .A(N111), .Y(n342) );
  INVX1_RVT U250 ( .A(A[11]), .Y(n117) );
  AO221X1_RVT U251 ( .A1(N176), .A2(n81), .A3(N252), .A4(n86), .A5(n261), .Y(
        n517) );
  AO221X1_RVT U252 ( .A1(N180), .A2(n81), .A3(N256), .A4(n86), .A5(n4), .Y(n45) );
  INVX1_RVT U253 ( .A(n9), .Y(n81) );
  INVX1_RVT U254 ( .A(n1), .Y(n86) );
  INVX0_RVT U255 ( .A(N179), .Y(n46) );
  OAI221X1_RVT U256 ( .A1(n46), .A2(n9), .A3(n47), .A4(n48), .A5(n49), .Y(n514) );
  AOI22X1_RVT U257 ( .A1(N204), .A2(n83), .A3(n103), .A4(n255), .Y(n49) );
  AOI221X1_RVT U258 ( .A1(N181), .A2(n81), .A3(N257), .A4(n86), .A5(n5), .Y(
        n50) );
  OAI221X1_RVT U259 ( .A1(N163), .A2(n324), .A3(N162), .A4(n326), .A5(n317), 
        .Y(n54) );
  INVX1_RVT U260 ( .A(n142), .Y(n139) );
  INVX1_RVT U261 ( .A(n155), .Y(n154) );
  INVX0_RVT U262 ( .A(\sub_1_root_add_170/carry[5] ), .Y(n145) );
  NAND2X0_RVT U263 ( .A1(n140), .A2(n145), .Y(n284) );
  NAND2X0_RVT U264 ( .A1(n146), .A2(n742), .Y(\sub_1_root_add_170/carry[7] )
         );
  AO21X1_RVT U265 ( .A1(B[22]), .A2(n142), .A3(n365), .Y(N516) );
  NAND2X0_RVT U266 ( .A1(next_state[0]), .A2(n144), .Y(n380) );
  NAND2X0_RVT U267 ( .A1(sel[0]), .A2(sel[1]), .Y(n608) );
  NAND2X0_RVT U268 ( .A1(n738), .A2(N516), .Y(n151) );
  AO21X1_RVT U269 ( .A1(n297), .A2(E[0]), .A3(n150), .Y(n149) );
  INVX0_RVT U270 ( .A(n558), .Y(n286) );
  AO22X1_RVT U271 ( .A1(E[0]), .A2(n286), .A3(N438), .A4(n519), .Y(n148) );
  AO221X1_RVT U272 ( .A1(n149), .A2(n289), .A3(N505), .A4(n513), .A5(n148), 
        .Y(n508) );
  NAND2X0_RVT U273 ( .A1(n150), .A2(n739), .Y(n155) );
  AO21X1_RVT U274 ( .A1(E[1]), .A2(n151), .A3(n154), .Y(n153) );
  AO22X1_RVT U275 ( .A1(n286), .A2(E[1]), .A3(N439), .A4(n519), .Y(n152) );
  AO221X1_RVT U276 ( .A1(n153), .A2(n289), .A3(N506), .A4(n513), .A5(n152), 
        .Y(n538) );
  NAND2X0_RVT U277 ( .A1(n154), .A2(n743), .Y(n159) );
  AO21X1_RVT U278 ( .A1(E[2]), .A2(n155), .A3(n158), .Y(n157) );
  AO22X1_RVT U279 ( .A1(n286), .A2(E[2]), .A3(N440), .A4(n519), .Y(n156) );
  AO221X1_RVT U280 ( .A1(n157), .A2(n289), .A3(N507), .A4(n513), .A5(n156), 
        .Y(n541) );
  NAND2X0_RVT U281 ( .A1(n158), .A2(n744), .Y(n163) );
  AO21X1_RVT U282 ( .A1(E[3]), .A2(n159), .A3(n162), .Y(n161) );
  AO22X1_RVT U283 ( .A1(n286), .A2(E[3]), .A3(N441), .A4(n519), .Y(n160) );
  AO221X1_RVT U284 ( .A1(n161), .A2(n289), .A3(N508), .A4(n513), .A5(n160), 
        .Y(n544) );
  NAND2X0_RVT U285 ( .A1(n162), .A2(n141), .Y(n167) );
  AO21X1_RVT U286 ( .A1(E[4]), .A2(n163), .A3(n166), .Y(n165) );
  AO22X1_RVT U287 ( .A1(n286), .A2(E[4]), .A3(N442), .A4(n519), .Y(n164) );
  AO221X1_RVT U288 ( .A1(n165), .A2(n289), .A3(N509), .A4(n513), .A5(n164), 
        .Y(n547) );
  NAND2X0_RVT U289 ( .A1(n166), .A2(n140), .Y(n171) );
  AO21X1_RVT U290 ( .A1(E[5]), .A2(n167), .A3(n170), .Y(n169) );
  AO22X1_RVT U291 ( .A1(n286), .A2(E[5]), .A3(N443), .A4(n519), .Y(n168) );
  AO221X1_RVT U292 ( .A1(n169), .A2(n289), .A3(N510), .A4(n513), .A5(n168), 
        .Y(n550) );
  NAND2X0_RVT U293 ( .A1(n170), .A2(n742), .Y(n277) );
  AO22X1_RVT U294 ( .A1(n286), .A2(E[6]), .A3(N444), .A4(n519), .Y(n172) );
  AO221X1_RVT U295 ( .A1(n173), .A2(n289), .A3(N511), .A4(n513), .A5(n172), 
        .Y(n553) );
  AO22X1_RVT U296 ( .A1(N500), .A2(n2), .A3(N359), .A4(n368), .Y(n554) );
  XOR2X1_RVT U297 ( .A1(E[7]), .A2(n174), .Y(n175) );
  AO22X1_RVT U298 ( .A1(n175), .A2(n289), .A3(n286), .A4(E[7]), .Y(n557) );
  INVX0_RVT U299 ( .A(n379), .Y(n292) );
  INVX0_RVT U300 ( .A(N167), .Y(n176) );
  AO221X1_RVT U301 ( .A1(N187), .A2(n81), .A3(N263), .A4(n85), .A5(n7), .Y(
        n506) );
  AO22X1_RVT U302 ( .A1(N211), .A2(n84), .A3(n104), .A4(n288), .Y(n177) );
  AO221X1_RVT U303 ( .A1(N186), .A2(n82), .A3(N262), .A4(n85), .A5(n177), .Y(
        n507) );
  AND3X1_RVT U304 ( .A1(n628), .A2(n635), .A3(n616), .Y(n178) );
  NAND3X0_RVT U305 ( .A1(n290), .A2(n292), .A3(n178), .Y(n280) );
  MUX21X1_RVT U306 ( .A1(div[46]), .A2(n139), .S0(n179), .Y(n423) );
  MUX21X1_RVT U307 ( .A1(div[45]), .A2(A[21]), .S0(n179), .Y(n422) );
  MUX21X1_RVT U308 ( .A1(div[44]), .A2(n136), .S0(n179), .Y(n421) );
  MUX21X1_RVT U309 ( .A1(div[43]), .A2(n132), .S0(n179), .Y(n420) );
  MUX21X1_RVT U310 ( .A1(div[42]), .A2(A[18]), .S0(n179), .Y(n419) );
  MUX21X1_RVT U311 ( .A1(div[41]), .A2(A[17]), .S0(n179), .Y(n418) );
  MUX21X1_RVT U312 ( .A1(div[40]), .A2(A[16]), .S0(n179), .Y(n417) );
  MUX21X1_RVT U313 ( .A1(div[39]), .A2(n122), .S0(n179), .Y(n416) );
  MUX21X1_RVT U314 ( .A1(div[38]), .A2(A[14]), .S0(n179), .Y(n415) );
  MUX21X1_RVT U315 ( .A1(div[37]), .A2(A[13]), .S0(n179), .Y(n414) );
  MUX21X1_RVT U316 ( .A1(div[36]), .A2(A[12]), .S0(n68), .Y(n413) );
  MUX21X1_RVT U317 ( .A1(div[35]), .A2(A[11]), .S0(n68), .Y(n412) );
  MUX21X1_RVT U318 ( .A1(div[34]), .A2(A[10]), .S0(n68), .Y(n411) );
  MUX21X1_RVT U319 ( .A1(div[33]), .A2(A[9]), .S0(n68), .Y(n410) );
  MUX21X1_RVT U320 ( .A1(div[32]), .A2(A[8]), .S0(n68), .Y(n409) );
  MUX21X1_RVT U321 ( .A1(div[31]), .A2(A[7]), .S0(n68), .Y(n408) );
  MUX21X1_RVT U322 ( .A1(div[30]), .A2(A[6]), .S0(n68), .Y(n407) );
  MUX21X1_RVT U323 ( .A1(div[29]), .A2(A[5]), .S0(n68), .Y(n406) );
  MUX21X1_RVT U324 ( .A1(div[28]), .A2(A[4]), .S0(n68), .Y(n405) );
  MUX21X1_RVT U325 ( .A1(div[27]), .A2(A[3]), .S0(n68), .Y(n404) );
  MUX21X1_RVT U326 ( .A1(div[26]), .A2(A[2]), .S0(n68), .Y(n403) );
  MUX21X1_RVT U327 ( .A1(div[25]), .A2(A[1]), .S0(n68), .Y(n402) );
  MUX21X1_RVT U328 ( .A1(div[24]), .A2(A[0]), .S0(n67), .Y(n401) );
  MUX21X1_RVT U329 ( .A1(divider[22]), .A2(B[22]), .S0(n67), .Y(n473) );
  MUX21X1_RVT U330 ( .A1(divider[21]), .A2(B[21]), .S0(n67), .Y(n474) );
  MUX21X1_RVT U331 ( .A1(divider[20]), .A2(B[20]), .S0(n67), .Y(n475) );
  MUX21X1_RVT U332 ( .A1(divider[19]), .A2(B[19]), .S0(n67), .Y(n476) );
  MUX21X1_RVT U333 ( .A1(divider[18]), .A2(B[18]), .S0(n67), .Y(n477) );
  MUX21X1_RVT U334 ( .A1(divider[17]), .A2(B[17]), .S0(n67), .Y(n478) );
  MUX21X1_RVT U335 ( .A1(divider[16]), .A2(B[16]), .S0(n67), .Y(n479) );
  MUX21X1_RVT U336 ( .A1(divider[15]), .A2(B[15]), .S0(n67), .Y(n480) );
  MUX21X1_RVT U337 ( .A1(divider[14]), .A2(B[14]), .S0(n67), .Y(n481) );
  MUX21X1_RVT U338 ( .A1(divider[13]), .A2(B[13]), .S0(n67), .Y(n482) );
  MUX21X1_RVT U339 ( .A1(divider[12]), .A2(B[12]), .S0(n67), .Y(n483) );
  MUX21X1_RVT U340 ( .A1(divider[11]), .A2(B[11]), .S0(n66), .Y(n484) );
  MUX21X1_RVT U341 ( .A1(divider[10]), .A2(B[10]), .S0(n66), .Y(n485) );
  MUX21X1_RVT U342 ( .A1(divider[9]), .A2(B[9]), .S0(n66), .Y(n486) );
  MUX21X1_RVT U343 ( .A1(divider[8]), .A2(B[8]), .S0(n66), .Y(n487) );
  MUX21X1_RVT U344 ( .A1(divider[7]), .A2(B[7]), .S0(n66), .Y(n488) );
  MUX21X1_RVT U345 ( .A1(divider[6]), .A2(B[6]), .S0(n66), .Y(n489) );
  MUX21X1_RVT U346 ( .A1(divider[5]), .A2(B[5]), .S0(n66), .Y(n490) );
  MUX21X1_RVT U347 ( .A1(divider[4]), .A2(B[4]), .S0(n66), .Y(n491) );
  MUX21X1_RVT U348 ( .A1(divider[3]), .A2(B[3]), .S0(n66), .Y(n492) );
  MUX21X1_RVT U349 ( .A1(divider[2]), .A2(B[2]), .S0(n66), .Y(n493) );
  MUX21X1_RVT U350 ( .A1(divider[1]), .A2(B[1]), .S0(n66), .Y(n494) );
  MUX21X1_RVT U351 ( .A1(divider[0]), .A2(B[0]), .S0(n66), .Y(n495) );
  AO222X1_RVT U352 ( .A1(N527), .A2(n41), .A3(N536), .A4(n10), .A5(
        quotient[23]), .A6(n574), .Y(n400) );
  AO222X1_RVT U353 ( .A1(N526), .A2(n41), .A3(N527), .A4(n10), .A5(
        quotient[22]), .A6(n574), .Y(n399) );
  AO222X1_RVT U354 ( .A1(N525), .A2(n41), .A3(N526), .A4(n10), .A5(
        quotient[21]), .A6(n574), .Y(n398) );
  AO222X1_RVT U355 ( .A1(N524), .A2(n41), .A3(N525), .A4(n10), .A5(
        quotient[20]), .A6(n574), .Y(n397) );
  AO222X1_RVT U356 ( .A1(N523), .A2(n41), .A3(N524), .A4(n10), .A5(
        quotient[19]), .A6(n574), .Y(n396) );
  AO222X1_RVT U357 ( .A1(N522), .A2(n41), .A3(N523), .A4(n10), .A5(
        quotient[18]), .A6(n574), .Y(n395) );
  AO222X1_RVT U358 ( .A1(N521), .A2(n41), .A3(N522), .A4(n10), .A5(
        quotient[17]), .A6(n574), .Y(n394) );
  AO222X1_RVT U359 ( .A1(N520), .A2(n41), .A3(N521), .A4(n10), .A5(
        quotient[16]), .A6(n574), .Y(n393) );
  AO222X1_RVT U360 ( .A1(quotient[15]), .A2(n574), .A3(N520), .A4(n10), .A5(
        n41), .A6(N519), .Y(n392) );
  NAND4X0_RVT U361 ( .A1(N641), .A2(quotient[16]), .A3(quotient[15]), .A4(n290), .Y(n591) );
  NAND3X0_RVT U362 ( .A1(n634), .A2(n42), .A3(n292), .Y(n281) );
  AO21X1_RVT U363 ( .A1(n568), .A2(n143), .A3(n180), .Y(n183) );
  NAND2X0_RVT U364 ( .A1(n183), .A2(n292), .Y(n181) );
  NAND2X0_RVT U365 ( .A1(n11), .A2(n183), .Y(n182) );
  AO222X1_RVT U366 ( .A1(N400), .A2(n78), .A3(n76), .A4(n287), .A5(n70), .A6(
        M1M2[39]), .Y(n433) );
  AO222X1_RVT U367 ( .A1(N401), .A2(n77), .A3(n76), .A4(M1M2[39]), .A5(n69), 
        .A6(M1M2[40]), .Y(n432) );
  AO222X1_RVT U368 ( .A1(N402), .A2(n77), .A3(n76), .A4(M1M2[40]), .A5(n69), 
        .A6(M1M2[41]), .Y(n431) );
  AO222X1_RVT U369 ( .A1(N403), .A2(n77), .A3(n76), .A4(M1M2[41]), .A5(n69), 
        .A6(M1M2[42]), .Y(n430) );
  AO222X1_RVT U370 ( .A1(N404), .A2(n77), .A3(n76), .A4(M1M2[42]), .A5(n69), 
        .A6(M1M2[43]), .Y(n429) );
  AO222X1_RVT U371 ( .A1(N405), .A2(n77), .A3(n76), .A4(M1M2[43]), .A5(n69), 
        .A6(M1M2[44]), .Y(n428) );
  AO222X1_RVT U372 ( .A1(N406), .A2(n77), .A3(n76), .A4(M1M2[44]), .A5(n69), 
        .A6(M1M2[45]), .Y(n427) );
  AO222X1_RVT U373 ( .A1(N407), .A2(n77), .A3(n76), .A4(M1M2[45]), .A5(n69), 
        .A6(M1M2[46]), .Y(n426) );
  AO222X1_RVT U374 ( .A1(N408), .A2(n77), .A3(n76), .A4(M1M2[46]), .A5(n69), 
        .A6(n279), .Y(n531) );
  AO22X1_RVT U375 ( .A1(N361), .A2(n80), .A3(n72), .A4(n184), .Y(n472) );
  AO222X1_RVT U376 ( .A1(N362), .A2(n77), .A3(n76), .A4(n184), .A5(n69), .A6(
        n185), .Y(n471) );
  AO222X1_RVT U377 ( .A1(N363), .A2(n77), .A3(n76), .A4(n185), .A5(n69), .A6(
        n186), .Y(n470) );
  AO222X1_RVT U378 ( .A1(N364), .A2(n77), .A3(n75), .A4(n186), .A5(n69), .A6(
        n187), .Y(n469) );
  AO222X1_RVT U379 ( .A1(N365), .A2(n78), .A3(n75), .A4(n187), .A5(n70), .A6(
        n188), .Y(n468) );
  AO222X1_RVT U380 ( .A1(N366), .A2(n78), .A3(n75), .A4(n188), .A5(n70), .A6(
        n189), .Y(n467) );
  AO222X1_RVT U381 ( .A1(N367), .A2(n78), .A3(n75), .A4(n189), .A5(n70), .A6(
        n190), .Y(n466) );
  AO222X1_RVT U382 ( .A1(N368), .A2(n78), .A3(n75), .A4(n190), .A5(n70), .A6(
        n191), .Y(n465) );
  AO222X1_RVT U383 ( .A1(N369), .A2(n78), .A3(n75), .A4(n191), .A5(n70), .A6(
        n192), .Y(n464) );
  AO222X1_RVT U384 ( .A1(N370), .A2(n78), .A3(n75), .A4(n192), .A5(n70), .A6(
        n193), .Y(n463) );
  AO222X1_RVT U385 ( .A1(N371), .A2(n78), .A3(n75), .A4(n193), .A5(n70), .A6(
        n194), .Y(n462) );
  AO222X1_RVT U386 ( .A1(N372), .A2(n78), .A3(n75), .A4(n194), .A5(n70), .A6(
        n195), .Y(n461) );
  AO222X1_RVT U387 ( .A1(N373), .A2(n78), .A3(n75), .A4(n195), .A5(n70), .A6(
        n196), .Y(n460) );
  AO222X1_RVT U388 ( .A1(N374), .A2(n78), .A3(n75), .A4(n196), .A5(n70), .A6(
        n197), .Y(n459) );
  AO222X1_RVT U389 ( .A1(N375), .A2(n78), .A3(n75), .A4(n197), .A5(n70), .A6(
        n198), .Y(n458) );
  AO222X1_RVT U390 ( .A1(N376), .A2(n79), .A3(n74), .A4(n198), .A5(n71), .A6(
        n199), .Y(n457) );
  AO222X1_RVT U391 ( .A1(N377), .A2(n79), .A3(n74), .A4(n199), .A5(n71), .A6(
        n200), .Y(n456) );
  AO222X1_RVT U392 ( .A1(N378), .A2(n79), .A3(n74), .A4(n200), .A5(n71), .A6(
        n201), .Y(n455) );
  AO222X1_RVT U393 ( .A1(N379), .A2(n79), .A3(n74), .A4(n201), .A5(n71), .A6(
        n203), .Y(n454) );
  AO222X1_RVT U394 ( .A1(N380), .A2(n79), .A3(n74), .A4(n203), .A5(n71), .A6(
        n204), .Y(n453) );
  AO222X1_RVT U395 ( .A1(N381), .A2(n79), .A3(n74), .A4(n204), .A5(n71), .A6(
        n205), .Y(n452) );
  AO222X1_RVT U396 ( .A1(N382), .A2(n79), .A3(n74), .A4(n205), .A5(n71), .A6(
        n206), .Y(n451) );
  AO222X1_RVT U397 ( .A1(N383), .A2(n79), .A3(n74), .A4(n206), .A5(n71), .A6(
        n207), .Y(n450) );
  AO222X1_RVT U398 ( .A1(N384), .A2(n79), .A3(n74), .A4(n207), .A5(n71), .A6(
        n208), .Y(n449) );
  AO222X1_RVT U399 ( .A1(N385), .A2(n79), .A3(n74), .A4(n208), .A5(n71), .A6(
        n209), .Y(n448) );
  AO222X1_RVT U400 ( .A1(N386), .A2(n79), .A3(n74), .A4(n209), .A5(n71), .A6(
        n210), .Y(n447) );
  AO222X1_RVT U401 ( .A1(N387), .A2(n79), .A3(n74), .A4(n210), .A5(n71), .A6(
        n212), .Y(n446) );
  AO222X1_RVT U402 ( .A1(N388), .A2(n80), .A3(n73), .A4(n212), .A5(n72), .A6(
        n213), .Y(n445) );
  AO222X1_RVT U403 ( .A1(N389), .A2(n80), .A3(n73), .A4(n213), .A5(n72), .A6(
        n215), .Y(n444) );
  AO222X1_RVT U404 ( .A1(N390), .A2(n80), .A3(n73), .A4(n215), .A5(n72), .A6(
        n216), .Y(n443) );
  AO222X1_RVT U405 ( .A1(N391), .A2(n80), .A3(n73), .A4(n216), .A5(n72), .A6(
        n218), .Y(n442) );
  AO222X1_RVT U406 ( .A1(N392), .A2(n80), .A3(n73), .A4(n218), .A5(n72), .A6(
        n219), .Y(n441) );
  AO222X1_RVT U407 ( .A1(N393), .A2(n80), .A3(n73), .A4(n219), .A5(n72), .A6(
        n221), .Y(n440) );
  AO222X1_RVT U408 ( .A1(N394), .A2(n80), .A3(n73), .A4(n221), .A5(n72), .A6(
        n222), .Y(n439) );
  AO222X1_RVT U409 ( .A1(N395), .A2(n80), .A3(n73), .A4(n222), .A5(n72), .A6(
        n224), .Y(n438) );
  AO222X1_RVT U410 ( .A1(N396), .A2(n80), .A3(n73), .A4(n224), .A5(n72), .A6(
        n225), .Y(n437) );
  AO222X1_RVT U411 ( .A1(N397), .A2(n80), .A3(n73), .A4(n225), .A5(n72), .A6(
        n227), .Y(n436) );
  AO222X1_RVT U412 ( .A1(N398), .A2(n80), .A3(n73), .A4(n227), .A5(n72), .A6(
        n228), .Y(n435) );
  AO222X1_RVT U413 ( .A1(N399), .A2(n77), .A3(n73), .A4(n228), .A5(n69), .A6(
        n287), .Y(n434) );
  AO22X1_RVT U414 ( .A1(N221), .A2(n84), .A3(n103), .A4(n229), .Y(n230) );
  AO22X1_RVT U415 ( .A1(N220), .A2(n84), .A3(n104), .A4(n231), .Y(n232) );
  AO221X1_RVT U416 ( .A1(N195), .A2(n82), .A3(N271), .A4(n85), .A5(n232), .Y(
        n498) );
  AO22X1_RVT U417 ( .A1(N219), .A2(n84), .A3(n104), .A4(n233), .Y(n234) );
  AO22X1_RVT U418 ( .A1(N218), .A2(n84), .A3(n104), .A4(n235), .Y(n236) );
  AO221X1_RVT U419 ( .A1(N193), .A2(n82), .A3(N269), .A4(n85), .A5(n236), .Y(
        n500) );
  AO22X1_RVT U420 ( .A1(N217), .A2(n84), .A3(n104), .A4(n237), .Y(n238) );
  AO221X1_RVT U421 ( .A1(N192), .A2(n82), .A3(N268), .A4(n85), .A5(n238), .Y(
        n501) );
  AO22X1_RVT U422 ( .A1(N216), .A2(n84), .A3(n104), .A4(n239), .Y(n240) );
  AO22X1_RVT U423 ( .A1(N215), .A2(n84), .A3(n104), .A4(n241), .Y(n242) );
  AO221X1_RVT U424 ( .A1(N190), .A2(n82), .A3(N266), .A4(n85), .A5(n242), .Y(
        n503) );
  AO22X1_RVT U425 ( .A1(N214), .A2(n84), .A3(n104), .A4(n243), .Y(n244) );
  AO221X1_RVT U426 ( .A1(N189), .A2(n82), .A3(N265), .A4(n85), .A5(n244), .Y(
        n504) );
  AO22X1_RVT U427 ( .A1(N213), .A2(n84), .A3(n104), .A4(n245), .Y(n246) );
  AO221X1_RVT U428 ( .A1(N188), .A2(n82), .A3(N264), .A4(n85), .A5(n246), .Y(
        n505) );
  AO22X1_RVT U429 ( .A1(N210), .A2(n84), .A3(n104), .A4(n247), .Y(n248) );
  AO22X1_RVT U430 ( .A1(N209), .A2(n84), .A3(n104), .A4(n249), .Y(n250) );
  AO22X1_RVT U431 ( .A1(N207), .A2(n83), .A3(n103), .A4(n252), .Y(n253) );
  AO221X1_RVT U432 ( .A1(N182), .A2(n81), .A3(N258), .A4(n86), .A5(n253), .Y(
        n511) );
  AO22X1_RVT U433 ( .A1(N203), .A2(n83), .A3(n103), .A4(n256), .Y(n257) );
  AO221X1_RVT U434 ( .A1(N178), .A2(n81), .A3(N254), .A4(n86), .A5(n257), .Y(
        n515) );
  AO22X1_RVT U435 ( .A1(N202), .A2(n83), .A3(n103), .A4(n258), .Y(n259) );
  AO221X1_RVT U436 ( .A1(N177), .A2(n81), .A3(N253), .A4(n86), .A5(n259), .Y(
        n516) );
  AO22X1_RVT U437 ( .A1(N201), .A2(n83), .A3(n104), .A4(n260), .Y(n261) );
  AO22X1_RVT U438 ( .A1(N200), .A2(n83), .A3(n103), .A4(n262), .Y(n263) );
  AO221X1_RVT U439 ( .A1(N175), .A2(n81), .A3(N251), .A4(n86), .A5(n263), .Y(
        n518) );
  AO22X1_RVT U440 ( .A1(N199), .A2(n83), .A3(n103), .A4(n264), .Y(n265) );
  AO22X1_RVT U441 ( .A1(N198), .A2(n83), .A3(n103), .A4(n266), .Y(n267) );
  AND3X1_RVT U442 ( .A1(n717), .A2(n721), .A3(n716), .Y(n269) );
  NAND4X0_RVT U443 ( .A1(n737), .A2(n736), .A3(n735), .A4(n269), .Y(n276) );
  AND4X1_RVT U444 ( .A1(n713), .A2(n715), .A3(n724), .A4(n723), .Y(n270) );
  NAND4X0_RVT U445 ( .A1(n720), .A2(n722), .A3(n718), .A4(n270), .Y(n275) );
  AND3X1_RVT U446 ( .A1(n719), .A2(n714), .A3(n732), .Y(n271) );
  NAND4X0_RVT U447 ( .A1(n727), .A2(n726), .A3(n725), .A4(n271), .Y(n274) );
  AND3X1_RVT U448 ( .A1(n730), .A2(n729), .A3(n731), .Y(n272) );
  NAND4X0_RVT U449 ( .A1(n734), .A2(n733), .A3(n728), .A4(n272), .Y(n273) );
  OR4X1_RVT U450 ( .A1(n276), .A2(n275), .A3(n274), .A4(n273), .Y(n610) );
  NAND4X0_RVT U451 ( .A1(n611), .A2(n376), .A3(n11), .A4(n610), .Y(n636) );
  NAND2X0_RVT U452 ( .A1(n568), .A2(n279), .Y(n637) );
  AND3X1_RVT U453 ( .A1(n281), .A2(n104), .A3(n280), .Y(n638) );
  NAND3X0_RVT U454 ( .A1(quotient[15]), .A2(quotient[16]), .A3(n587), .Y(n697)
         );
  AO22X1_RVT U455 ( .A1(N634), .A2(n20), .A3(n39), .A4(quotient[16]), .Y(n689)
         );
  AO22X1_RVT U456 ( .A1(N635), .A2(n20), .A3(quotient[17]), .A4(n39), .Y(n690)
         );
  AO22X1_RVT U457 ( .A1(N636), .A2(n20), .A3(quotient[18]), .A4(n39), .Y(n691)
         );
  AO22X1_RVT U458 ( .A1(N637), .A2(n20), .A3(quotient[19]), .A4(n39), .Y(n692)
         );
  AO22X1_RVT U459 ( .A1(N638), .A2(n20), .A3(quotient[20]), .A4(n39), .Y(n693)
         );
  AO22X1_RVT U460 ( .A1(N639), .A2(n20), .A3(quotient[21]), .A4(n39), .Y(n694)
         );
  NAND4X0_RVT U461 ( .A1(E[6]), .A2(E[7]), .A3(E[0]), .A4(E[1]), .Y(n702) );
  NAND4X0_RVT U462 ( .A1(E[4]), .A2(E[5]), .A3(E[2]), .A4(E[3]), .Y(n703) );
  XOR2X1_RVT U463 ( .A1(E[7]), .A2(n283), .Y(N491) );
  AO21X1_RVT U464 ( .A1(E[6]), .A2(n284), .A3(n283), .Y(N490) );
  AOI222X1_RVT U465 ( .A1(N501), .A2(n2), .A3(n286), .A4(n285), .A5(N360), 
        .A6(n368), .Y(n745) );
  XNOR2X1_RVT U466 ( .A1(\sub_1_root_sub_0_root_sub_122/carry[7] ), .A2(N437), 
        .Y(N350) );
  AND2X1_RVT U467 ( .A1(B[29]), .A2(\sub_1_root_sub_0_root_sub_122/carry[6] ), 
        .Y(\sub_1_root_sub_0_root_sub_122/carry[7] ) );
  XOR2X1_RVT U468 ( .A1(B[29]), .A2(\sub_1_root_sub_0_root_sub_122/carry[6] ), 
        .Y(N349) );
  AND2X1_RVT U469 ( .A1(B[28]), .A2(\sub_1_root_sub_0_root_sub_122/carry[5] ), 
        .Y(\sub_1_root_sub_0_root_sub_122/carry[6] ) );
  XOR2X1_RVT U470 ( .A1(B[28]), .A2(\sub_1_root_sub_0_root_sub_122/carry[5] ), 
        .Y(N348) );
  AND2X1_RVT U471 ( .A1(B[27]), .A2(\sub_1_root_sub_0_root_sub_122/carry[4] ), 
        .Y(\sub_1_root_sub_0_root_sub_122/carry[5] ) );
  XOR2X1_RVT U472 ( .A1(B[27]), .A2(\sub_1_root_sub_0_root_sub_122/carry[4] ), 
        .Y(N347) );
  AND2X1_RVT U473 ( .A1(B[26]), .A2(\sub_1_root_sub_0_root_sub_122/carry[3] ), 
        .Y(\sub_1_root_sub_0_root_sub_122/carry[4] ) );
  XOR2X1_RVT U474 ( .A1(B[26]), .A2(\sub_1_root_sub_0_root_sub_122/carry[3] ), 
        .Y(N346) );
  AND2X1_RVT U475 ( .A1(B[25]), .A2(\sub_1_root_sub_0_root_sub_122/carry[2] ), 
        .Y(\sub_1_root_sub_0_root_sub_122/carry[3] ) );
  XOR2X1_RVT U476 ( .A1(B[25]), .A2(\sub_1_root_sub_0_root_sub_122/carry[2] ), 
        .Y(N345) );
  AND2X1_RVT U477 ( .A1(B[24]), .A2(n31), .Y(
        \sub_1_root_sub_0_root_sub_122/carry[2] ) );
  XOR2X1_RVT U478 ( .A1(B[24]), .A2(n32), .Y(N344) );
  XNOR2X1_RVT U479 ( .A1(n285), .A2(\sub_1_root_add_170/carry[8] ), .Y(N492)
         );
  OR2X1_RVT U480 ( .A1(E[7]), .A2(\sub_1_root_add_170/carry[7] ), .Y(
        \sub_1_root_add_170/carry[8] ) );
  XNOR2X1_RVT U481 ( .A1(\sub_1_root_add_170/carry[5] ), .A2(E[5]), .Y(N489)
         );
  OR2X1_RVT U482 ( .A1(E[0]), .A2(n105), .Y(\sub_1_root_add_170/carry[1] ) );
  XNOR2X1_RVT U483 ( .A1(n105), .A2(E[0]), .Y(N484) );
  XNOR2X1_RVT U484 ( .A1(N437), .A2(\sub_143/carry[7] ), .Y(N424) );
  AND2X1_RVT U485 ( .A1(B[29]), .A2(\sub_143/carry[6] ), .Y(\sub_143/carry[7] ) );
  XOR2X1_RVT U486 ( .A1(B[29]), .A2(\sub_143/carry[6] ), .Y(N423) );
  AND2X1_RVT U487 ( .A1(B[28]), .A2(\sub_143/carry[5] ), .Y(\sub_143/carry[6] ) );
  XOR2X1_RVT U488 ( .A1(B[28]), .A2(\sub_143/carry[5] ), .Y(N422) );
  AND2X1_RVT U489 ( .A1(B[27]), .A2(\sub_143/carry[4] ), .Y(\sub_143/carry[5] ) );
  XOR2X1_RVT U490 ( .A1(B[27]), .A2(\sub_143/carry[4] ), .Y(N421) );
  AND2X1_RVT U491 ( .A1(B[26]), .A2(\sub_143/carry[3] ), .Y(\sub_143/carry[4] ) );
  XOR2X1_RVT U492 ( .A1(B[26]), .A2(\sub_143/carry[3] ), .Y(N420) );
  AND2X1_RVT U493 ( .A1(B[25]), .A2(\sub_143/carry[2] ), .Y(\sub_143/carry[3] ) );
  XOR2X1_RVT U494 ( .A1(B[25]), .A2(\sub_143/carry[2] ), .Y(N419) );
  AND2X1_RVT U495 ( .A1(B[24]), .A2(n31), .Y(\sub_143/carry[2] ) );
  XOR2X1_RVT U496 ( .A1(B[24]), .A2(n31), .Y(N418) );
  AND2X1_RVT U497 ( .A1(N143), .A2(n342), .Y(n298) );
  AND2X1_RVT U498 ( .A1(n298), .A2(n321), .Y(n299) );
  OA222X1_RVT U499 ( .A1(N145), .A2(n320), .A3(N144), .A4(n299), .A5(n298), 
        .A6(n321), .Y(n300) );
  AO221X1_RVT U500 ( .A1(N145), .A2(n320), .A3(N146), .A4(n319), .A5(n300), 
        .Y(n301) );
  OA221X1_RVT U501 ( .A1(N147), .A2(n336), .A3(N146), .A4(n319), .A5(n301), 
        .Y(n302) );
  AO221X1_RVT U504 ( .A1(N147), .A2(n336), .A3(N148), .A4(n335), .A5(n302), 
        .Y(n303) );
  OA221X1_RVT U505 ( .A1(N149), .A2(n334), .A3(N148), .A4(n335), .A5(n303), 
        .Y(n304) );
  AO221X1_RVT U506 ( .A1(N149), .A2(n334), .A3(N150), .A4(n333), .A5(n304), 
        .Y(n305) );
  OA221X1_RVT U507 ( .A1(N151), .A2(n331), .A3(N150), .A4(n333), .A5(n305), 
        .Y(n306) );
  OA221X1_RVT U508 ( .A1(N152), .A2(n330), .A3(N153), .A4(n341), .A5(n307), 
        .Y(n308) );
  AO221X1_RVT U509 ( .A1(N153), .A2(n341), .A3(N154), .A4(n340), .A5(n308), 
        .Y(n309) );
  OA221X1_RVT U510 ( .A1(N155), .A2(n339), .A3(N154), .A4(n340), .A5(n309), 
        .Y(n310) );
  AO221X1_RVT U511 ( .A1(N155), .A2(n339), .A3(N156), .A4(n338), .A5(n310), 
        .Y(n311) );
  OA221X1_RVT U512 ( .A1(N157), .A2(n332), .A3(N156), .A4(n338), .A5(n311), 
        .Y(n312) );
  AO221X1_RVT U513 ( .A1(N157), .A2(n332), .A3(N158), .A4(n337), .A5(n312), 
        .Y(n313) );
  OA221X1_RVT U514 ( .A1(N159), .A2(n329), .A3(N158), .A4(n337), .A5(n313), 
        .Y(n314) );
  OA221X1_RVT U515 ( .A1(N161), .A2(n327), .A3(N160), .A4(n328), .A5(n315), 
        .Y(n316) );
  AO221X1_RVT U516 ( .A1(N161), .A2(n327), .A3(N162), .A4(n326), .A5(n316), 
        .Y(n317) );
  OA221X1_RVT U517 ( .A1(N165), .A2(n325), .A3(N164), .A4(n322), .A5(n37), .Y(
        n318) );
  AND2X1_RVT U518 ( .A1(B[0]), .A2(n106), .Y(n343) );
  AND2X1_RVT U519 ( .A1(n343), .A2(n107), .Y(n344) );
  OA222X1_RVT U520 ( .A1(B[2]), .A2(n108), .A3(B[1]), .A4(n344), .A5(n343), 
        .A6(n107), .Y(n345) );
  AO221X1_RVT U521 ( .A1(B[2]), .A2(n108), .A3(B[3]), .A4(n109), .A5(n345), 
        .Y(n346) );
  OA221X1_RVT U522 ( .A1(B[4]), .A2(n110), .A3(B[3]), .A4(n109), .A5(n346), 
        .Y(n347) );
  AO221X1_RVT U523 ( .A1(B[4]), .A2(n110), .A3(B[5]), .A4(n111), .A5(n347), 
        .Y(n348) );
  OA221X1_RVT U524 ( .A1(B[6]), .A2(n112), .A3(B[5]), .A4(n111), .A5(n348), 
        .Y(n349) );
  AO221X1_RVT U525 ( .A1(B[6]), .A2(n112), .A3(B[7]), .A4(n113), .A5(n349), 
        .Y(n350) );
  OA221X1_RVT U526 ( .A1(B[8]), .A2(n114), .A3(B[7]), .A4(n113), .A5(n350), 
        .Y(n351) );
  AO221X1_RVT U527 ( .A1(B[8]), .A2(n114), .A3(B[9]), .A4(n115), .A5(n351), 
        .Y(n352) );
  OA221X1_RVT U528 ( .A1(B[9]), .A2(n115), .A3(B[10]), .A4(n116), .A5(n352), 
        .Y(n353) );
  AO221X1_RVT U529 ( .A1(B[10]), .A2(n116), .A3(B[11]), .A4(n117), .A5(n353), 
        .Y(n354) );
  OA221X1_RVT U530 ( .A1(B[12]), .A2(n118), .A3(B[11]), .A4(n117), .A5(n354), 
        .Y(n355) );
  AO221X1_RVT U531 ( .A1(B[12]), .A2(n118), .A3(B[13]), .A4(n119), .A5(n355), 
        .Y(n356) );
  OA221X1_RVT U532 ( .A1(B[14]), .A2(n120), .A3(B[13]), .A4(n119), .A5(n356), 
        .Y(n357) );
  AO221X1_RVT U533 ( .A1(B[14]), .A2(n120), .A3(B[15]), .A4(n124), .A5(n357), 
        .Y(n358) );
  OA221X1_RVT U534 ( .A1(B[16]), .A2(n126), .A3(B[15]), .A4(n124), .A5(n358), 
        .Y(n359) );
  AO221X1_RVT U535 ( .A1(B[16]), .A2(n126), .A3(B[17]), .A4(n128), .A5(n359), 
        .Y(n360) );
  OA221X1_RVT U536 ( .A1(B[18]), .A2(n130), .A3(B[17]), .A4(n128), .A5(n360), 
        .Y(n361) );
  AO221X1_RVT U537 ( .A1(B[18]), .A2(n130), .A3(B[19]), .A4(n134), .A5(n361), 
        .Y(n362) );
  OA221X1_RVT U538 ( .A1(B[20]), .A2(n137), .A3(B[19]), .A4(n134), .A5(n362), 
        .Y(n363) );
  AO221X1_RVT U539 ( .A1(B[20]), .A2(n137), .A3(B[21]), .A4(n138), .A5(n363), 
        .Y(n364) );
  OA221X1_RVT U540 ( .A1(B[22]), .A2(n142), .A3(B[21]), .A4(n138), .A5(n364), 
        .Y(n365) );
  AND4X1_RVT U541 ( .A1(N333), .A2(N332), .A3(N336), .A4(N335), .Y(n366) );
  AND4X1_RVT U542 ( .A1(N330), .A2(N334), .A3(N331), .A4(n366), .Y(n367) );
  AOI222X1_RVT U543 ( .A1(n369), .A2(Y[21]), .A3(result[21]), .A4(n370), .A5(
        N579), .A6(n371), .Y(n746) );
  AOI222X1_RVT U544 ( .A1(n369), .A2(Y[20]), .A3(result[20]), .A4(n370), .A5(
        N578), .A6(n371), .Y(n747) );
  AOI222X1_RVT U545 ( .A1(n369), .A2(Y[19]), .A3(result[19]), .A4(n370), .A5(
        N577), .A6(n371), .Y(n748) );
  AOI222X1_RVT U546 ( .A1(n369), .A2(Y[18]), .A3(result[18]), .A4(n370), .A5(
        N576), .A6(n371), .Y(n749) );
  AOI222X1_RVT U547 ( .A1(n369), .A2(Y[17]), .A3(result[17]), .A4(n370), .A5(
        N575), .A6(n371), .Y(n750) );
  AOI222X1_RVT U548 ( .A1(n369), .A2(Y[16]), .A3(result[16]), .A4(n370), .A5(
        N574), .A6(n371), .Y(n751) );
  AOI222X1_RVT U549 ( .A1(n369), .A2(Y[15]), .A3(result[15]), .A4(n370), .A5(
        N573), .A6(n371), .Y(n752) );
  NOR4X0_RVT U550 ( .A1(n372), .A2(n373), .A3(n374), .A4(sel[1]), .Y(n371) );
  AND3X1_RVT U551 ( .A1(n375), .A2(n376), .A3(n377), .Y(n370) );
  NAND2X0_RVT U552 ( .A1(n378), .A2(n379), .Y(n532) );
  MUX21X1_RVT U553 ( .A1(n380), .A2(n381), .S0(n11), .Y(n378) );
  OR3X1_RVT U554 ( .A1(n499), .A2(n502), .A3(n508), .Y(n530) );
  AO22X1_RVT U555 ( .A1(n521), .A2(A[23]), .A3(n535), .A4(n32), .Y(n502) );
  AO22X1_RVT U556 ( .A1(N352), .A2(n368), .A3(N493), .A4(n2), .Y(n499) );
  OR3X1_RVT U557 ( .A1(n536), .A2(n537), .A3(n538), .Y(n529) );
  AO22X1_RVT U558 ( .A1(n521), .A2(A[24]), .A3(n535), .A4(B[24]), .Y(n537) );
  AO22X1_RVT U559 ( .A1(N353), .A2(n368), .A3(N494), .A4(n2), .Y(n536) );
  OR3X1_RVT U560 ( .A1(n539), .A2(n540), .A3(n541), .Y(n528) );
  AO22X1_RVT U561 ( .A1(n521), .A2(A[25]), .A3(n535), .A4(B[25]), .Y(n540) );
  AO22X1_RVT U562 ( .A1(N354), .A2(n368), .A3(N495), .A4(n2), .Y(n539) );
  OR3X1_RVT U563 ( .A1(n542), .A2(n543), .A3(n544), .Y(n527) );
  AO22X1_RVT U564 ( .A1(n521), .A2(A[26]), .A3(n535), .A4(B[26]), .Y(n543) );
  AO22X1_RVT U565 ( .A1(N355), .A2(n368), .A3(N496), .A4(n2), .Y(n542) );
  OR3X1_RVT U566 ( .A1(n545), .A2(n546), .A3(n547), .Y(n526) );
  AO22X1_RVT U567 ( .A1(n521), .A2(A[27]), .A3(n535), .A4(B[27]), .Y(n546) );
  AO22X1_RVT U568 ( .A1(N356), .A2(n368), .A3(N497), .A4(n2), .Y(n545) );
  OR3X1_RVT U569 ( .A1(n548), .A2(n549), .A3(n550), .Y(n525) );
  AO22X1_RVT U570 ( .A1(n521), .A2(A[28]), .A3(n535), .A4(B[28]), .Y(n549) );
  AO22X1_RVT U571 ( .A1(N357), .A2(n368), .A3(N498), .A4(n2), .Y(n548) );
  OR3X1_RVT U572 ( .A1(n551), .A2(n552), .A3(n553), .Y(n524) );
  AO22X1_RVT U573 ( .A1(n521), .A2(A[29]), .A3(n535), .A4(B[29]), .Y(n552) );
  AO22X1_RVT U574 ( .A1(N358), .A2(n368), .A3(N499), .A4(n2), .Y(n551) );
  OR3X1_RVT U575 ( .A1(n554), .A2(n555), .A3(n556), .Y(n523) );
  AO221X1_RVT U576 ( .A1(N512), .A2(n513), .A3(N445), .A4(n519), .A5(n557), 
        .Y(n556) );
  AO22X1_RVT U577 ( .A1(n521), .A2(n65), .A3(n535), .A4(N437), .Y(n555) );
  AND3X1_RVT U578 ( .A1(n559), .A2(n376), .A3(n97), .Y(n535) );
  AND3X1_RVT U579 ( .A1(n95), .A2(n376), .A3(n559), .Y(n521) );
  MUX21X1_RVT U580 ( .A1(n562), .A2(n144), .S0(n379), .Y(n522) );
  AO21X1_RVT U581 ( .A1(n103), .A2(n564), .A3(n565), .Y(n496) );
  MUX21X1_RVT U582 ( .A1(n85), .A2(n566), .S0(A[31]), .Y(n565) );
  AO21X1_RVT U583 ( .A1(N167), .A2(n40), .A3(n83), .Y(n566) );
  AO22X1_RVT U584 ( .A1(error), .A2(n144), .A3(n292), .A4(n569), .Y(n425) );
  MUX21X1_RVT U585 ( .A1(n570), .A2(over_flow), .S0(n571), .Y(n424) );
  OA221X1_RVT U586 ( .A1(n572), .A2(n373), .A3(n573), .A4(n379), .A5(n144), 
        .Y(n571) );
  NAND2X0_RVT U587 ( .A1(n373), .A2(n379), .Y(n570) );
  MUX21X1_RVT U588 ( .A1(Y[22]), .A2(n575), .S0(n576), .Y(n391) );
  AO22X1_RVT U589 ( .A1(n577), .A2(n578), .A3(n579), .A4(n580), .Y(n575) );
  AND2X1_RVT U590 ( .A1(n581), .A2(n291), .Y(n579) );
  NAND4X0_RVT U591 ( .A1(n582), .A2(n583), .A3(n584), .A4(n585), .Y(n578) );
  NAND3X0_RVT U592 ( .A1(n586), .A2(n587), .A3(n572), .Y(n585) );
  NAND2X0_RVT U593 ( .A1(n588), .A2(n589), .Y(n586) );
  NAND4X0_RVT U594 ( .A1(N580), .A2(M_sum[15]), .A3(n288), .A4(n376), .Y(n589)
         );
  AO21X1_RVT U595 ( .A1(n590), .A2(n591), .A3(n592), .Y(n588) );
  INVX0_RVT U596 ( .A(n593), .Y(n592) );
  NAND4X0_RVT U597 ( .A1(N611), .A2(n561), .A3(n287), .A4(M1M2[39]), .Y(n590)
         );
  NAND3X0_RVT U598 ( .A1(n377), .A2(n376), .A3(result[22]), .Y(n584) );
  AND2X1_RVT U599 ( .A1(n572), .A2(n372), .Y(n377) );
  NAND3X0_RVT U600 ( .A1(n288), .A2(n587), .A3(M_sum[15]), .Y(n372) );
  NAND3X0_RVT U601 ( .A1(quotient[23]), .A2(n290), .A3(n594), .Y(n583) );
  NAND3X0_RVT U602 ( .A1(n561), .A2(M1M2[46]), .A3(n595), .Y(n582) );
  AO221X1_RVT U603 ( .A1(n596), .A2(E[0]), .A3(n369), .A4(Y[23]), .A5(n597), 
        .Y(n390) );
  AO221X1_RVT U604 ( .A1(n596), .A2(E[1]), .A3(n369), .A4(Y[24]), .A5(n597), 
        .Y(n389) );
  AO221X1_RVT U605 ( .A1(n596), .A2(E[2]), .A3(n369), .A4(Y[25]), .A5(n597), 
        .Y(n388) );
  AO221X1_RVT U606 ( .A1(n596), .A2(E[3]), .A3(n369), .A4(Y[26]), .A5(n597), 
        .Y(n387) );
  AO221X1_RVT U607 ( .A1(n596), .A2(E[4]), .A3(n369), .A4(Y[27]), .A5(n597), 
        .Y(n386) );
  AO221X1_RVT U608 ( .A1(n596), .A2(E[5]), .A3(n369), .A4(Y[28]), .A5(n597), 
        .Y(n385) );
  AO221X1_RVT U609 ( .A1(n596), .A2(E[6]), .A3(n369), .A4(Y[29]), .A5(n597), 
        .Y(n384) );
  AO221X1_RVT U610 ( .A1(n596), .A2(E[7]), .A3(n369), .A4(Y[30]), .A5(n597), 
        .Y(n383) );
  AO21X1_RVT U611 ( .A1(n596), .A2(n374), .A3(n598), .Y(n597) );
  AND4X1_RVT U612 ( .A1(n599), .A2(n576), .A3(n581), .A4(n291), .Y(n598) );
  NAND2X0_RVT U613 ( .A1(n600), .A2(n573), .Y(n599) );
  INVX0_RVT U614 ( .A(n580), .Y(n600) );
  NAND2X0_RVT U615 ( .A1(n601), .A2(sel[1]), .Y(n580) );
  INVX0_RVT U616 ( .A(n572), .Y(n374) );
  AO221X1_RVT U617 ( .A1(n602), .A2(n603), .A3(n369), .A4(Y[31]), .A5(n604), 
        .Y(n382) );
  AND3X1_RVT U618 ( .A1(n564), .A2(n376), .A3(n596), .Y(n604) );
  AO22X1_RVT U619 ( .A1(n605), .A2(n576), .A3(n596), .A4(n606), .Y(n603) );
  NAND2X0_RVT U620 ( .A1(n607), .A2(n608), .Y(n606) );
  AO221X1_RVT U621 ( .A1(n292), .A2(n562), .A3(n609), .A4(n11), .A5(n375), .Y(
        n576) );
  INVX0_RVT U622 ( .A(n381), .Y(n609) );
  AO21X1_RVT U623 ( .A1(n610), .A2(n611), .A3(sel[1]), .Y(n381) );
  NAND3X0_RVT U624 ( .A1(n612), .A2(n613), .A3(n614), .Y(n562) );
  OA22X1_RVT U625 ( .A1(n615), .A2(n42), .A3(n616), .A4(n608), .Y(n614) );
  INVX0_RVT U626 ( .A(n569), .Y(n612) );
  NAND2X0_RVT U627 ( .A1(n601), .A2(n617), .Y(n569) );
  NAND3X0_RVT U628 ( .A1(n563), .A2(n376), .A3(n618), .Y(n617) );
  AOI22X1_RVT U629 ( .A1(n561), .A2(n619), .A3(n290), .A4(n620), .Y(n601) );
  AO21X1_RVT U630 ( .A1(n621), .A2(n622), .A3(n618), .Y(n620) );
  NAND3X0_RVT U631 ( .A1(n623), .A2(n615), .A3(n613), .Y(n605) );
  AND2X1_RVT U632 ( .A1(n573), .A2(n624), .Y(n613) );
  NAND3X0_RVT U633 ( .A1(n561), .A2(n625), .A3(n626), .Y(n624) );
  NAND2X0_RVT U634 ( .A1(n627), .A2(n628), .Y(n625) );
  AND2X1_RVT U635 ( .A1(n629), .A2(n630), .Y(n573) );
  NAND3X0_RVT U636 ( .A1(n561), .A2(n631), .A3(n626), .Y(n630) );
  AO22X1_RVT U637 ( .A1(n621), .A2(n632), .A3(n622), .A4(n633), .Y(n619) );
  NAND3X0_RVT U638 ( .A1(n290), .A2(n627), .A3(n621), .Y(n629) );
  INVX0_RVT U639 ( .A(n634), .Y(n615) );
  NAND3X0_RVT U640 ( .A1(n628), .A2(n635), .A3(n290), .Y(n623) );
  AO222X1_RVT U641 ( .A1(N446), .A2(n519), .A3(N513), .A4(n513), .A5(N545), 
        .A6(n289), .Y(n323) );
  AND2X1_RVT U642 ( .A1(n292), .A2(n558), .Y(n559) );
  NAND4X0_RVT U643 ( .A1(n636), .A2(n574), .A3(n637), .A4(n638), .Y(n558) );
  AOI22X1_RVT U644 ( .A1(N424), .A2(n64), .A3(n639), .A4(n640), .Y(n616) );
  OR2X1_RVT U645 ( .A1(n64), .A2(N424), .Y(n640) );
  AO21X1_RVT U646 ( .A1(N423), .A2(n63), .A3(n641), .Y(n639) );
  OA221X1_RVT U647 ( .A1(N422), .A2(n62), .A3(N423), .A4(n63), .A5(n642), .Y(
        n641) );
  AO221X1_RVT U648 ( .A1(N421), .A2(n643), .A3(N422), .A4(n62), .A5(n644), .Y(
        n642) );
  OA221X1_RVT U649 ( .A1(N420), .A2(n61), .A3(N421), .A4(n643), .A5(n645), .Y(
        n644) );
  AO222X1_RVT U650 ( .A1(n646), .A2(n60), .A3(N419), .A4(n647), .A5(N420), 
        .A6(n61), .Y(n645) );
  OR2X1_RVT U651 ( .A1(n60), .A2(n646), .Y(n647) );
  OA22X1_RVT U652 ( .A1(n648), .A2(n649), .A3(N418), .A4(n650), .Y(n646) );
  AO21X1_RVT U653 ( .A1(N418), .A2(n650), .A3(n55), .Y(n649) );
  INVX0_RVT U654 ( .A(n628), .Y(n621) );
  OR2X1_RVT U655 ( .A1(n651), .A2(n652), .Y(n628) );
  NAND4X0_RVT U656 ( .A1(n55), .A2(n653), .A3(n56), .A4(n57), .Y(n652) );
  NAND4X0_RVT U657 ( .A1(n58), .A2(n654), .A3(n59), .A4(n655), .Y(n651) );
  INVX0_RVT U658 ( .A(n627), .Y(n622) );
  OR2X1_RVT U659 ( .A1(n656), .A2(n657), .Y(n627) );
  NAND4X0_RVT U660 ( .A1(n648), .A2(n650), .A3(n60), .A4(n61), .Y(n657) );
  NAND4X0_RVT U661 ( .A1(n643), .A2(n62), .A3(n63), .A4(n64), .Y(n656) );
  INVX0_RVT U662 ( .A(A[27]), .Y(n643) );
  NAND2X0_RVT U663 ( .A1(n658), .A2(n659), .Y(n631) );
  NAND2X0_RVT U664 ( .A1(n618), .A2(n563), .Y(n660) );
  INVX0_RVT U665 ( .A(n567), .Y(n563) );
  XOR2X1_RVT U666 ( .A1(n661), .A2(n602), .Y(n567) );
  XOR2X1_RVT U667 ( .A1(A[31]), .A2(B[31]), .Y(n602) );
  INVX0_RVT U668 ( .A(n635), .Y(n618) );
  NAND2X0_RVT U669 ( .A1(n632), .A2(n633), .Y(n635) );
  INVX0_RVT U670 ( .A(n659), .Y(n633) );
  NAND4X0_RVT U671 ( .A1(n662), .A2(n663), .A3(n664), .A4(n665), .Y(n659) );
  NOR4X0_RVT U672 ( .A1(n666), .A2(n667), .A3(n668), .A4(n669), .Y(n665) );
  OR4X1_RVT U673 ( .A1(B[16]), .A2(B[17]), .A3(B[18]), .A4(B[19]), .Y(n669) );
  OR4X1_RVT U674 ( .A1(B[1]), .A2(B[20]), .A3(B[21]), .A4(B[22]), .Y(n668) );
  OR4X1_RVT U675 ( .A1(B[2]), .A2(B[3]), .A3(B[4]), .A4(B[5]), .Y(n667) );
  OR4X1_RVT U676 ( .A1(B[6]), .A2(B[7]), .A3(B[8]), .A4(B[9]), .Y(n666) );
  AND4X1_RVT U677 ( .A1(B[29]), .A2(B[28]), .A3(N437), .A4(n670), .Y(n664) );
  AND4X1_RVT U678 ( .A1(B[27]), .A2(B[26]), .A3(B[25]), .A4(B[24]), .Y(n670)
         );
  NOR4X0_RVT U679 ( .A1(B[12]), .A2(B[13]), .A3(B[14]), .A4(B[15]), .Y(n663)
         );
  NOR4X0_RVT U680 ( .A1(n55), .A2(B[0]), .A3(B[10]), .A4(B[11]), .Y(n662) );
  INVX0_RVT U681 ( .A(n658), .Y(n632) );
  NAND4X0_RVT U682 ( .A1(n671), .A2(n672), .A3(n673), .A4(n674), .Y(n658) );
  NOR4X0_RVT U683 ( .A1(n675), .A2(n676), .A3(n677), .A4(n678), .Y(n674) );
  OR4X1_RVT U684 ( .A1(A[16]), .A2(A[17]), .A3(A[18]), .A4(n132), .Y(n678) );
  OR4X1_RVT U685 ( .A1(A[1]), .A2(n136), .A3(A[21]), .A4(n139), .Y(n677) );
  OR4X1_RVT U686 ( .A1(A[2]), .A2(A[3]), .A3(A[4]), .A4(A[5]), .Y(n676) );
  OR4X1_RVT U687 ( .A1(A[6]), .A2(A[7]), .A3(A[8]), .A4(A[9]), .Y(n675) );
  AND4X1_RVT U688 ( .A1(A[29]), .A2(A[28]), .A3(n65), .A4(n679), .Y(n673) );
  NOR4X0_RVT U689 ( .A1(A[12]), .A2(A[13]), .A3(A[14]), .A4(n122), .Y(n672) );
  NOR4X0_RVT U690 ( .A1(n648), .A2(A[0]), .A3(A[10]), .A4(A[11]), .Y(n671) );
  AND2X1_RVT U691 ( .A1(n11), .A2(n561), .Y(n568) );
  INVX0_RVT U692 ( .A(sel[1]), .Y(n376) );
  NAND4X0_RVT U693 ( .A1(n140), .A2(n680), .A3(n742), .A4(n681), .Y(n611) );
  AND2X1_RVT U694 ( .A1(n740), .A2(n741), .Y(n681) );
  AO21X1_RVT U695 ( .A1(shifted[4]), .A2(n141), .A3(n682), .Y(n680) );
  OA221X1_RVT U696 ( .A1(shifted[3]), .A2(n744), .A3(shifted[4]), .A4(n141), 
        .A5(n683), .Y(n682) );
  AO221X1_RVT U697 ( .A1(shifted[2]), .A2(n743), .A3(shifted[3]), .A4(n744), 
        .A5(n684), .Y(n683) );
  OA222X1_RVT U698 ( .A1(shifted[2]), .A2(n743), .A3(shifted[1]), .A4(n685), 
        .A5(n739), .A6(n686), .Y(n684) );
  AND2X1_RVT U699 ( .A1(n739), .A2(n686), .Y(n685) );
  AND2X1_RVT U700 ( .A1(shifted[0]), .A2(n738), .Y(n686) );
  NAND3X0_RVT U701 ( .A1(n291), .A2(n144), .A3(n581), .Y(n379) );
  AO221X1_RVT U702 ( .A1(N604), .A2(n687), .A3(n688), .A4(M1M2[39]), .A5(n689), 
        .Y(n226) );
  AO221X1_RVT U703 ( .A1(N605), .A2(n687), .A3(n688), .A4(M1M2[40]), .A5(n690), 
        .Y(n223) );
  AO221X1_RVT U704 ( .A1(N606), .A2(n687), .A3(n688), .A4(M1M2[41]), .A5(n691), 
        .Y(n220) );
  AO221X1_RVT U705 ( .A1(N607), .A2(n687), .A3(n688), .A4(M1M2[42]), .A5(n692), 
        .Y(n217) );
  AO221X1_RVT U706 ( .A1(N608), .A2(n687), .A3(n688), .A4(M1M2[43]), .A5(n693), 
        .Y(n214) );
  AO221X1_RVT U707 ( .A1(N609), .A2(n687), .A3(n688), .A4(M1M2[44]), .A5(n694), 
        .Y(n211) );
  AO221X1_RVT U708 ( .A1(N610), .A2(n687), .A3(n688), .A4(M1M2[45]), .A5(n695), 
        .Y(n202) );
  AO22X1_RVT U709 ( .A1(N640), .A2(n20), .A3(n39), .A4(quotient[22]), .Y(n695)
         );
  AND2X1_RVT U710 ( .A1(n696), .A2(n697), .Y(n594) );
  AND3X1_RVT U711 ( .A1(n375), .A2(n561), .A3(n595), .Y(n688) );
  AND2X1_RVT U712 ( .A1(n696), .A2(n698), .Y(n595) );
  AND4X1_RVT U713 ( .A1(n699), .A2(n696), .A3(n375), .A4(n561), .Y(n687) );
  NAND2X0_RVT U714 ( .A1(sel[1]), .A2(n661), .Y(n607) );
  INVX0_RVT U715 ( .A(sel[0]), .Y(n661) );
  INVX0_RVT U716 ( .A(n373), .Y(n375) );
  NAND2X0_RVT U717 ( .A1(n577), .A2(n144), .Y(n373) );
  AND2X1_RVT U718 ( .A1(next_state[1]), .A2(n581), .Y(n577) );
  AND2X1_RVT U719 ( .A1(n572), .A2(n593), .Y(n696) );
  OR2X1_RVT U720 ( .A1(n700), .A2(n701), .Y(n593) );
  NAND4X0_RVT U721 ( .A1(n740), .A2(n742), .A3(n140), .A4(n141), .Y(n701) );
  NAND4X0_RVT U722 ( .A1(n744), .A2(n743), .A3(n739), .A4(n738), .Y(n700) );
  OA21X1_RVT U723 ( .A1(n702), .A2(n703), .A3(n741), .Y(n572) );
  INVX0_RVT U724 ( .A(n698), .Y(n699) );
  NAND3X0_RVT U725 ( .A1(M1M2[39]), .A2(n587), .A3(n287), .Y(n698) );
  INVX0_RVT U726 ( .A(round_mode), .Y(n587) );
  OR2X1_RVT U727 ( .A1(N110), .A2(n94), .Y(N166) );
  MUX21X1_RVT U728 ( .A1(N109), .A2(n139), .S0(n93), .Y(N165) );
  MUX21X1_RVT U729 ( .A1(N108), .A2(A[21]), .S0(n93), .Y(N164) );
  MUX21X1_RVT U730 ( .A1(N107), .A2(n136), .S0(n93), .Y(N163) );
  MUX21X1_RVT U731 ( .A1(N106), .A2(n132), .S0(n93), .Y(N162) );
  MUX21X1_RVT U732 ( .A1(N105), .A2(A[18]), .S0(n93), .Y(N161) );
  MUX21X1_RVT U733 ( .A1(N104), .A2(A[17]), .S0(n93), .Y(N160) );
  MUX21X1_RVT U734 ( .A1(N103), .A2(A[16]), .S0(n93), .Y(N159) );
  MUX21X1_RVT U735 ( .A1(N101), .A2(A[14]), .S0(n92), .Y(N157) );
  MUX21X1_RVT U736 ( .A1(N100), .A2(A[13]), .S0(n92), .Y(N156) );
  MUX21X1_RVT U737 ( .A1(N98), .A2(A[11]), .S0(n90), .Y(N154) );
  MUX21X1_RVT U738 ( .A1(N97), .A2(A[10]), .S0(n90), .Y(N153) );
  MUX21X1_RVT U739 ( .A1(N96), .A2(A[9]), .S0(n89), .Y(N152) );
  MUX21X1_RVT U740 ( .A1(N93), .A2(A[6]), .S0(n92), .Y(N149) );
  MUX21X1_RVT U741 ( .A1(N92), .A2(A[5]), .S0(n88), .Y(N148) );
  MUX21X1_RVT U742 ( .A1(N91), .A2(A[4]), .S0(n91), .Y(N147) );
  MUX21X1_RVT U743 ( .A1(N89), .A2(A[2]), .S0(n87), .Y(N145) );
  MUX21X1_RVT U744 ( .A1(N88), .A2(A[1]), .S0(n87), .Y(N144) );
  OR2X1_RVT U745 ( .A1(n97), .A2(N78), .Y(N134) );
  MUX21X1_RVT U746 ( .A1(N77), .A2(B[22]), .S0(n101), .Y(N133) );
  MUX21X1_RVT U747 ( .A1(N76), .A2(B[21]), .S0(n101), .Y(N132) );
  MUX21X1_RVT U748 ( .A1(N75), .A2(B[20]), .S0(n101), .Y(N131) );
  MUX21X1_RVT U749 ( .A1(N74), .A2(B[19]), .S0(n102), .Y(N130) );
  MUX21X1_RVT U750 ( .A1(N73), .A2(B[18]), .S0(n101), .Y(N129) );
  MUX21X1_RVT U751 ( .A1(N72), .A2(B[17]), .S0(n101), .Y(N128) );
  MUX21X1_RVT U752 ( .A1(N71), .A2(B[16]), .S0(n101), .Y(N127) );
  MUX21X1_RVT U753 ( .A1(N70), .A2(B[15]), .S0(n101), .Y(N126) );
  MUX21X1_RVT U754 ( .A1(N69), .A2(B[14]), .S0(n101), .Y(N125) );
  MUX21X1_RVT U755 ( .A1(N68), .A2(B[13]), .S0(n101), .Y(N124) );
  MUX21X1_RVT U756 ( .A1(N67), .A2(B[12]), .S0(n101), .Y(N123) );
  MUX21X1_RVT U757 ( .A1(N66), .A2(B[11]), .S0(n102), .Y(N122) );
  MUX21X1_RVT U758 ( .A1(N65), .A2(B[10]), .S0(n102), .Y(N121) );
  MUX21X1_RVT U759 ( .A1(N64), .A2(B[9]), .S0(n102), .Y(N120) );
  MUX21X1_RVT U760 ( .A1(N63), .A2(B[8]), .S0(n102), .Y(N119) );
  MUX21X1_RVT U761 ( .A1(N62), .A2(B[7]), .S0(n102), .Y(N118) );
  MUX21X1_RVT U762 ( .A1(N61), .A2(B[6]), .S0(n102), .Y(N117) );
  MUX21X1_RVT U763 ( .A1(N60), .A2(B[5]), .S0(n102), .Y(N116) );
  MUX21X1_RVT U764 ( .A1(N59), .A2(B[4]), .S0(n102), .Y(N115) );
  MUX21X1_RVT U765 ( .A1(N58), .A2(B[3]), .S0(n102), .Y(N114) );
  MUX21X1_RVT U766 ( .A1(N57), .A2(B[2]), .S0(n102), .Y(N113) );
  MUX21X1_RVT U767 ( .A1(N56), .A2(B[1]), .S0(n102), .Y(N112) );
  MUX21X1_RVT U768 ( .A1(N55), .A2(B[0]), .S0(n101), .Y(N111) );
  AO22X1_RVT U769 ( .A1(n65), .A2(n655), .A3(n704), .A4(n705), .Y(n560) );
  NAND2X0_RVT U770 ( .A1(N437), .A2(n64), .Y(n705) );
  AO21X1_RVT U771 ( .A1(A[29]), .A2(n59), .A3(n706), .Y(n704) );
  OA221X1_RVT U772 ( .A1(A[28]), .A2(n654), .A3(A[29]), .A4(n59), .A5(n707), 
        .Y(n706) );
  AO221X1_RVT U773 ( .A1(A[27]), .A2(n58), .A3(A[28]), .A4(n654), .A5(n708), 
        .Y(n707) );
  OA221X1_RVT U774 ( .A1(A[26]), .A2(n57), .A3(A[27]), .A4(n58), .A5(n709), 
        .Y(n708) );
  AO222X1_RVT U775 ( .A1(A[25]), .A2(n710), .A3(n711), .A4(n56), .A5(A[26]), 
        .A6(n57), .Y(n709) );
  OR2X1_RVT U776 ( .A1(n710), .A2(A[25]), .Y(n711) );
  AO22X1_RVT U777 ( .A1(A[24]), .A2(n653), .A3(n712), .A4(A[23]), .Y(n710) );
  INVX0_RVT U778 ( .A(B[24]), .Y(n653) );
  INVX0_RVT U779 ( .A(B[28]), .Y(n654) );
  INVX0_RVT U780 ( .A(N437), .Y(n655) );
endmodule


module FPU ( clk, reset, A, B, sel, round_mode, start, error, over_flow, Y );
  input [31:0] A;
  input [31:0] B;
  input [1:0] sel;
  output [31:0] Y;
  input clk, reset, round_mode, start;
  output error, over_flow;
  wire   round_fpu, error_fpu, over_flow_fpu, n1, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128;
  wire   [31:0] A_fpu;
  wire   [31:0] B_fpu;
  wire   [1:0] sel_fpu;
  wire   [31:0] Y_fpu;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14;
  assign Y[14] = 1'b0;
  assign Y[13] = 1'b0;
  assign Y[12] = 1'b0;
  assign Y[11] = 1'b0;
  assign Y[10] = 1'b0;
  assign Y[9] = 1'b0;
  assign Y[8] = 1'b0;
  assign Y[7] = 1'b0;
  assign Y[6] = 1'b0;
  assign Y[5] = 1'b0;
  assign Y[4] = 1'b0;
  assign Y[3] = 1'b0;
  assign Y[2] = 1'b0;
  assign Y[1] = 1'b0;
  assign Y[0] = 1'b0;

  NAND2X0_RVT U5 ( .A1(reset), .A2(n119), .Y(n1) );
  FPU_CAL fpu_cal ( .clk(clk), .start(n112), .A({A_fpu[31:23], n105, 
        A_fpu[21:0]}), .B(B_fpu), .sel(sel_fpu), .round_mode(round_fpu), 
        .error(error_fpu), .over_flow(over_flow_fpu), .Y({Y_fpu[31:15], 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14}) );
  DFFARX1_RVT \A_fpu_reg[21]  ( .D(n94), .CLK(clk), .RSTB(n120), .Q(A_fpu[21])
         );
  DFFARX1_RVT \A_fpu_reg[22]  ( .D(n95), .CLK(clk), .RSTB(n120), .Q(n105) );
  DFFARX1_RVT \A_fpu_reg[10]  ( .D(n83), .CLK(clk), .RSTB(n121), .Q(A_fpu[10])
         );
  DFFARX1_RVT \B_fpu_reg[23]  ( .D(n64), .CLK(clk), .RSTB(n123), .Q(B_fpu[23])
         );
  DFFARX1_RVT \A_fpu_reg[23]  ( .D(n96), .CLK(clk), .RSTB(n120), .Q(A_fpu[23])
         );
  DFFX1_RVT over_flow_reg ( .D(n5), .CLK(clk), .Q(over_flow) );
  DFFX1_RVT error_reg ( .D(n4), .CLK(clk), .Q(error) );
  DFFARX1_RVT \Y_reg[15]  ( .D(n22), .CLK(clk), .RSTB(reset), .Q(Y[15]) );
  DFFARX1_RVT \Y_reg[16]  ( .D(n21), .CLK(clk), .RSTB(reset), .Q(Y[16]) );
  DFFARX1_RVT \Y_reg[17]  ( .D(n20), .CLK(clk), .RSTB(n126), .Q(Y[17]) );
  DFFARX1_RVT \Y_reg[18]  ( .D(n19), .CLK(clk), .RSTB(n126), .Q(Y[18]) );
  DFFARX1_RVT \Y_reg[19]  ( .D(n18), .CLK(clk), .RSTB(n126), .Q(Y[19]) );
  DFFARX1_RVT \Y_reg[20]  ( .D(n17), .CLK(clk), .RSTB(n126), .Q(Y[20]) );
  DFFARX1_RVT \Y_reg[21]  ( .D(n16), .CLK(clk), .RSTB(n126), .Q(Y[21]) );
  DFFARX1_RVT \Y_reg[22]  ( .D(n15), .CLK(clk), .RSTB(n126), .Q(Y[22]) );
  DFFARX1_RVT \Y_reg[23]  ( .D(n14), .CLK(clk), .RSTB(n126), .Q(Y[23]) );
  DFFARX1_RVT \Y_reg[24]  ( .D(n13), .CLK(clk), .RSTB(n126), .Q(Y[24]) );
  DFFARX1_RVT \Y_reg[25]  ( .D(n12), .CLK(clk), .RSTB(n126), .Q(Y[25]) );
  DFFARX1_RVT \Y_reg[26]  ( .D(n11), .CLK(clk), .RSTB(n126), .Q(Y[26]) );
  DFFARX1_RVT \Y_reg[27]  ( .D(n10), .CLK(clk), .RSTB(n126), .Q(Y[27]) );
  DFFARX1_RVT \Y_reg[28]  ( .D(n9), .CLK(clk), .RSTB(n126), .Q(Y[28]) );
  DFFARX1_RVT \Y_reg[29]  ( .D(n8), .CLK(clk), .RSTB(reset), .Q(Y[29]) );
  DFFARX1_RVT \Y_reg[30]  ( .D(n7), .CLK(clk), .RSTB(reset), .Q(Y[30]) );
  DFFARX1_RVT \Y_reg[31]  ( .D(n6), .CLK(clk), .RSTB(reset), .Q(Y[31]) );
  DFFARX1_RVT round_fpu_reg ( .D(n38), .CLK(clk), .RSTB(n125), .Q(round_fpu)
         );
  DFFARX1_RVT \A_fpu_reg[1]  ( .D(n74), .CLK(clk), .RSTB(n122), .Q(A_fpu[1])
         );
  DFFARX1_RVT \A_fpu_reg[2]  ( .D(n75), .CLK(clk), .RSTB(n122), .Q(A_fpu[2])
         );
  DFFARX1_RVT \A_fpu_reg[4]  ( .D(n77), .CLK(clk), .RSTB(n122), .Q(A_fpu[4])
         );
  DFFARX1_RVT \A_fpu_reg[3]  ( .D(n76), .CLK(clk), .RSTB(n122), .Q(A_fpu[3])
         );
  DFFARX1_RVT \A_fpu_reg[5]  ( .D(n78), .CLK(clk), .RSTB(n122), .Q(A_fpu[5])
         );
  DFFARX1_RVT \A_fpu_reg[0]  ( .D(n73), .CLK(clk), .RSTB(n122), .Q(A_fpu[0])
         );
  DFFARX1_RVT \A_fpu_reg[6]  ( .D(n79), .CLK(clk), .RSTB(n122), .Q(A_fpu[6])
         );
  DFFARX1_RVT \A_fpu_reg[7]  ( .D(n80), .CLK(clk), .RSTB(n122), .Q(A_fpu[7])
         );
  DFFARX1_RVT \A_fpu_reg[20]  ( .D(n93), .CLK(clk), .RSTB(n120), .Q(A_fpu[20])
         );
  DFFARX1_RVT \A_fpu_reg[18]  ( .D(n91), .CLK(clk), .RSTB(n121), .Q(A_fpu[18])
         );
  DFFARX1_RVT \A_fpu_reg[19]  ( .D(n92), .CLK(clk), .RSTB(n121), .Q(A_fpu[19])
         );
  DFFARX1_RVT \A_fpu_reg[16]  ( .D(n89), .CLK(clk), .RSTB(n121), .Q(A_fpu[16])
         );
  DFFARX1_RVT \A_fpu_reg[17]  ( .D(n90), .CLK(clk), .RSTB(n121), .Q(A_fpu[17])
         );
  DFFARX1_RVT \A_fpu_reg[14]  ( .D(n87), .CLK(clk), .RSTB(n121), .Q(A_fpu[14])
         );
  DFFARX1_RVT \A_fpu_reg[15]  ( .D(n88), .CLK(clk), .RSTB(n121), .Q(A_fpu[15])
         );
  DFFARX1_RVT \A_fpu_reg[13]  ( .D(n86), .CLK(clk), .RSTB(n121), .Q(A_fpu[13])
         );
  DFFARX1_RVT \A_fpu_reg[12]  ( .D(n85), .CLK(clk), .RSTB(n121), .Q(A_fpu[12])
         );
  DFFARX1_RVT \A_fpu_reg[9]  ( .D(n82), .CLK(clk), .RSTB(n121), .Q(A_fpu[9])
         );
  DFFARX1_RVT \A_fpu_reg[8]  ( .D(n81), .CLK(clk), .RSTB(n121), .Q(A_fpu[8])
         );
  DFFARX1_RVT \B_fpu_reg[31]  ( .D(n72), .CLK(clk), .RSTB(n122), .Q(B_fpu[31])
         );
  DFFARX1_RVT \sel_fpu_reg[0]  ( .D(n39), .CLK(clk), .RSTB(n125), .Q(
        sel_fpu[0]) );
  DFFARX1_RVT \A_fpu_reg[31]  ( .D(n104), .CLK(clk), .RSTB(n120), .Q(A_fpu[31]) );
  DFFARX1_RVT \sel_fpu_reg[1]  ( .D(n40), .CLK(clk), .RSTB(n125), .Q(
        sel_fpu[1]) );
  DFFARX1_RVT \B_fpu_reg[0]  ( .D(n41), .CLK(clk), .RSTB(n125), .Q(B_fpu[0])
         );
  DFFARX1_RVT \B_fpu_reg[1]  ( .D(n42), .CLK(clk), .RSTB(n125), .Q(B_fpu[1])
         );
  DFFARX1_RVT \B_fpu_reg[2]  ( .D(n43), .CLK(clk), .RSTB(n125), .Q(B_fpu[2])
         );
  DFFARX1_RVT \B_fpu_reg[20]  ( .D(n61), .CLK(clk), .RSTB(n123), .Q(B_fpu[20])
         );
  DFFARX1_RVT \B_fpu_reg[6]  ( .D(n47), .CLK(clk), .RSTB(n124), .Q(B_fpu[6])
         );
  DFFARX1_RVT \B_fpu_reg[16]  ( .D(n57), .CLK(clk), .RSTB(n123), .Q(B_fpu[16])
         );
  DFFARX1_RVT \B_fpu_reg[27]  ( .D(n68), .CLK(clk), .RSTB(n123), .Q(B_fpu[27])
         );
  DFFARX1_RVT \A_fpu_reg[27]  ( .D(n100), .CLK(clk), .RSTB(n120), .Q(A_fpu[27]) );
  DFFARX1_RVT \B_fpu_reg[26]  ( .D(n67), .CLK(clk), .RSTB(n123), .Q(B_fpu[26])
         );
  DFFARX1_RVT \A_fpu_reg[26]  ( .D(n99), .CLK(clk), .RSTB(n120), .Q(A_fpu[26])
         );
  DFFARX1_RVT \B_fpu_reg[28]  ( .D(n69), .CLK(clk), .RSTB(n122), .Q(B_fpu[28])
         );
  DFFARX1_RVT \B_fpu_reg[29]  ( .D(n70), .CLK(clk), .RSTB(n122), .Q(B_fpu[29])
         );
  DFFARX1_RVT \A_fpu_reg[28]  ( .D(n101), .CLK(clk), .RSTB(n120), .Q(A_fpu[28]) );
  DFFARX1_RVT \A_fpu_reg[29]  ( .D(n102), .CLK(clk), .RSTB(n120), .Q(A_fpu[29]) );
  DFFARX1_RVT \B_fpu_reg[25]  ( .D(n66), .CLK(clk), .RSTB(n123), .Q(B_fpu[25])
         );
  DFFARX1_RVT \A_fpu_reg[25]  ( .D(n98), .CLK(clk), .RSTB(n120), .Q(A_fpu[25])
         );
  DFFARX1_RVT \B_fpu_reg[30]  ( .D(n71), .CLK(clk), .RSTB(n122), .Q(B_fpu[30])
         );
  DFFARX1_RVT \A_fpu_reg[30]  ( .D(n103), .CLK(clk), .RSTB(n120), .Q(A_fpu[30]) );
  DFFARX1_RVT \B_fpu_reg[12]  ( .D(n53), .CLK(clk), .RSTB(n124), .Q(B_fpu[12])
         );
  DFFARX1_RVT \B_fpu_reg[4]  ( .D(n45), .CLK(clk), .RSTB(n124), .Q(B_fpu[4])
         );
  DFFARX1_RVT \B_fpu_reg[8]  ( .D(n49), .CLK(clk), .RSTB(n124), .Q(B_fpu[8])
         );
  DFFARX1_RVT \B_fpu_reg[9]  ( .D(n50), .CLK(clk), .RSTB(n124), .Q(B_fpu[9])
         );
  DFFARX1_RVT \B_fpu_reg[14]  ( .D(n55), .CLK(clk), .RSTB(n124), .Q(B_fpu[14])
         );
  DFFARX1_RVT \B_fpu_reg[22]  ( .D(n63), .CLK(clk), .RSTB(n123), .Q(B_fpu[22])
         );
  DFFARX1_RVT \B_fpu_reg[3]  ( .D(n44), .CLK(clk), .RSTB(n125), .Q(B_fpu[3])
         );
  DFFARX1_RVT \B_fpu_reg[17]  ( .D(n58), .CLK(clk), .RSTB(n123), .Q(B_fpu[17])
         );
  DFFARX1_RVT \B_fpu_reg[7]  ( .D(n48), .CLK(clk), .RSTB(n124), .Q(B_fpu[7])
         );
  DFFARX1_RVT \B_fpu_reg[13]  ( .D(n54), .CLK(clk), .RSTB(n124), .Q(B_fpu[13])
         );
  DFFARX1_RVT \B_fpu_reg[18]  ( .D(n59), .CLK(clk), .RSTB(n123), .Q(B_fpu[18])
         );
  DFFARX1_RVT \B_fpu_reg[21]  ( .D(n62), .CLK(clk), .RSTB(n123), .Q(B_fpu[21])
         );
  DFFARX1_RVT \B_fpu_reg[5]  ( .D(n46), .CLK(clk), .RSTB(n124), .Q(B_fpu[5])
         );
  DFFARX1_RVT \B_fpu_reg[10]  ( .D(n51), .CLK(clk), .RSTB(n124), .Q(B_fpu[10])
         );
  DFFARX1_RVT \B_fpu_reg[11]  ( .D(n52), .CLK(clk), .RSTB(n124), .Q(B_fpu[11])
         );
  DFFARX1_RVT \B_fpu_reg[15]  ( .D(n56), .CLK(clk), .RSTB(n124), .Q(B_fpu[15])
         );
  DFFARX1_RVT \B_fpu_reg[19]  ( .D(n60), .CLK(clk), .RSTB(n123), .Q(B_fpu[19])
         );
  DFFARX1_RVT \B_fpu_reg[24]  ( .D(n65), .CLK(clk), .RSTB(n123), .Q(B_fpu[24])
         );
  DFFARX1_RVT \A_fpu_reg[24]  ( .D(n97), .CLK(clk), .RSTB(n120), .Q(A_fpu[24])
         );
  DFFARX1_RVT \A_fpu_reg[11]  ( .D(n84), .CLK(clk), .RSTB(n121), .Q(A_fpu[11])
         );
  INVX1_RVT U106 ( .A(n1), .Y(n128) );
  INVX1_RVT U107 ( .A(n127), .Y(n120) );
  INVX1_RVT U108 ( .A(n127), .Y(n123) );
  INVX1_RVT U109 ( .A(n127), .Y(n121) );
  INVX1_RVT U110 ( .A(n127), .Y(n126) );
  INVX1_RVT U111 ( .A(n127), .Y(n124) );
  INVX1_RVT U112 ( .A(n127), .Y(n122) );
  INVX1_RVT U113 ( .A(n127), .Y(n125) );
  INVX1_RVT U114 ( .A(n113), .Y(n107) );
  INVX1_RVT U115 ( .A(n113), .Y(n108) );
  INVX1_RVT U116 ( .A(n113), .Y(n106) );
  INVX1_RVT U117 ( .A(n113), .Y(n112) );
  INVX1_RVT U118 ( .A(n113), .Y(n111) );
  INVX1_RVT U119 ( .A(n113), .Y(n109) );
  INVX1_RVT U120 ( .A(n113), .Y(n110) );
  AO22X1_RVT U121 ( .A1(n1), .A2(error), .A3(error_fpu), .A4(n128), .Y(n4) );
  AO22X1_RVT U122 ( .A1(over_flow), .A2(n1), .A3(over_flow_fpu), .A4(n128), 
        .Y(n5) );
  AO22X1_RVT U123 ( .A1(A_fpu[23]), .A2(n119), .A3(A[23]), .A4(n106), .Y(n96)
         );
  AO22X1_RVT U124 ( .A1(B_fpu[19]), .A2(n116), .A3(B[19]), .A4(n109), .Y(n60)
         );
  AO22X1_RVT U125 ( .A1(B_fpu[11]), .A2(n115), .A3(B[11]), .A4(n110), .Y(n52)
         );
  AO22X1_RVT U126 ( .A1(B_fpu[15]), .A2(n116), .A3(B[15]), .A4(n109), .Y(n56)
         );
  AO22X1_RVT U127 ( .A1(B_fpu[21]), .A2(n116), .A3(B[21]), .A4(n109), .Y(n62)
         );
  AO22X1_RVT U128 ( .A1(B_fpu[5]), .A2(n115), .A3(B[5]), .A4(n110), .Y(n46) );
  AO22X1_RVT U129 ( .A1(B_fpu[10]), .A2(n115), .A3(B[10]), .A4(n110), .Y(n51)
         );
  AO22X1_RVT U130 ( .A1(B_fpu[18]), .A2(n116), .A3(B[18]), .A4(n109), .Y(n59)
         );
  AO22X1_RVT U131 ( .A1(B_fpu[22]), .A2(n116), .A3(B[22]), .A4(n109), .Y(n63)
         );
  AO22X1_RVT U132 ( .A1(B_fpu[9]), .A2(n115), .A3(B[9]), .A4(n110), .Y(n50) );
  AO22X1_RVT U133 ( .A1(B_fpu[13]), .A2(n116), .A3(B[13]), .A4(n110), .Y(n54)
         );
  AO22X1_RVT U134 ( .A1(B_fpu[14]), .A2(n116), .A3(B[14]), .A4(n110), .Y(n55)
         );
  AO22X1_RVT U135 ( .A1(B_fpu[3]), .A2(n115), .A3(B[3]), .A4(n110), .Y(n44) );
  AO22X1_RVT U136 ( .A1(B_fpu[7]), .A2(n115), .A3(B[7]), .A4(n110), .Y(n48) );
  AO22X1_RVT U137 ( .A1(B_fpu[17]), .A2(n116), .A3(B[17]), .A4(n109), .Y(n58)
         );
  AO22X1_RVT U138 ( .A1(B_fpu[4]), .A2(n115), .A3(B[4]), .A4(n110), .Y(n45) );
  AO22X1_RVT U139 ( .A1(B_fpu[8]), .A2(n115), .A3(B[8]), .A4(n110), .Y(n49) );
  AO22X1_RVT U140 ( .A1(B_fpu[24]), .A2(n116), .A3(B[24]), .A4(n109), .Y(n65)
         );
  AO22X1_RVT U141 ( .A1(B_fpu[25]), .A2(n116), .A3(B[25]), .A4(n109), .Y(n66)
         );
  AO22X1_RVT U142 ( .A1(B_fpu[26]), .A2(n117), .A3(B[26]), .A4(n109), .Y(n67)
         );
  AO22X1_RVT U143 ( .A1(B_fpu[27]), .A2(n117), .A3(B[27]), .A4(n108), .Y(n68)
         );
  AO22X1_RVT U144 ( .A1(B_fpu[28]), .A2(n117), .A3(B[28]), .A4(n108), .Y(n69)
         );
  AO22X1_RVT U145 ( .A1(B_fpu[29]), .A2(n117), .A3(B[29]), .A4(n108), .Y(n70)
         );
  AO22X1_RVT U146 ( .A1(B_fpu[30]), .A2(n117), .A3(B[30]), .A4(n108), .Y(n71)
         );
  AO22X1_RVT U147 ( .A1(A_fpu[24]), .A2(n119), .A3(A[24]), .A4(n106), .Y(n97)
         );
  AO22X1_RVT U148 ( .A1(A_fpu[25]), .A2(n119), .A3(A[25]), .A4(n106), .Y(n98)
         );
  AO22X1_RVT U149 ( .A1(A_fpu[26]), .A2(n119), .A3(A[26]), .A4(n106), .Y(n99)
         );
  AO22X1_RVT U150 ( .A1(A_fpu[27]), .A2(n119), .A3(A[27]), .A4(n106), .Y(n100)
         );
  AO22X1_RVT U151 ( .A1(A_fpu[28]), .A2(n119), .A3(A[28]), .A4(n106), .Y(n101)
         );
  AO22X1_RVT U152 ( .A1(A_fpu[29]), .A2(n119), .A3(A[29]), .A4(n106), .Y(n102)
         );
  AO22X1_RVT U153 ( .A1(A_fpu[30]), .A2(n119), .A3(A[30]), .A4(n106), .Y(n103)
         );
  AO22X1_RVT U154 ( .A1(B_fpu[12]), .A2(n116), .A3(B[12]), .A4(n110), .Y(n53)
         );
  AO22X1_RVT U155 ( .A1(B_fpu[20]), .A2(n116), .A3(B[20]), .A4(n109), .Y(n61)
         );
  AO22X1_RVT U156 ( .A1(B_fpu[6]), .A2(n115), .A3(B[6]), .A4(n110), .Y(n47) );
  AO22X1_RVT U157 ( .A1(B_fpu[16]), .A2(n116), .A3(B[16]), .A4(n109), .Y(n57)
         );
  AO22X1_RVT U158 ( .A1(A_fpu[11]), .A2(n118), .A3(A[11]), .A4(n107), .Y(n84)
         );
  AO22X1_RVT U159 ( .A1(B_fpu[2]), .A2(n115), .A3(B[2]), .A4(n110), .Y(n43) );
  AO22X1_RVT U160 ( .A1(B_fpu[1]), .A2(n115), .A3(B[1]), .A4(n111), .Y(n42) );
  AO22X1_RVT U161 ( .A1(B_fpu[0]), .A2(n115), .A3(B[0]), .A4(n111), .Y(n41) );
  AO22X1_RVT U162 ( .A1(sel_fpu[1]), .A2(n115), .A3(sel[1]), .A4(n111), .Y(n40) );
  AO22X1_RVT U163 ( .A1(n112), .A2(Y[31]), .A3(Y_fpu[31]), .A4(n113), .Y(n6)
         );
  AO22X1_RVT U164 ( .A1(n112), .A2(Y[30]), .A3(Y_fpu[30]), .A4(n113), .Y(n7)
         );
  AO22X1_RVT U165 ( .A1(n112), .A2(Y[29]), .A3(Y_fpu[29]), .A4(n113), .Y(n8)
         );
  AO22X1_RVT U166 ( .A1(n112), .A2(Y[28]), .A3(Y_fpu[28]), .A4(n113), .Y(n9)
         );
  AO22X1_RVT U167 ( .A1(n112), .A2(Y[27]), .A3(Y_fpu[27]), .A4(n113), .Y(n10)
         );
  AO22X1_RVT U168 ( .A1(n112), .A2(Y[26]), .A3(Y_fpu[26]), .A4(n114), .Y(n11)
         );
  AO22X1_RVT U169 ( .A1(n112), .A2(Y[25]), .A3(Y_fpu[25]), .A4(n114), .Y(n12)
         );
  AO22X1_RVT U170 ( .A1(n112), .A2(Y[24]), .A3(Y_fpu[24]), .A4(n114), .Y(n13)
         );
  AO22X1_RVT U171 ( .A1(A_fpu[31]), .A2(n119), .A3(A[31]), .A4(n109), .Y(n104)
         );
  AO22X1_RVT U172 ( .A1(sel_fpu[0]), .A2(n115), .A3(sel[0]), .A4(n111), .Y(n39) );
  AO22X1_RVT U173 ( .A1(B_fpu[31]), .A2(n117), .A3(B[31]), .A4(n108), .Y(n72)
         );
  AO22X1_RVT U174 ( .A1(A_fpu[0]), .A2(n117), .A3(A[0]), .A4(n108), .Y(n73) );
  AO22X1_RVT U175 ( .A1(A_fpu[1]), .A2(n117), .A3(A[1]), .A4(n108), .Y(n74) );
  AO22X1_RVT U176 ( .A1(A_fpu[2]), .A2(n117), .A3(A[2]), .A4(n108), .Y(n75) );
  AO22X1_RVT U177 ( .A1(A_fpu[3]), .A2(n117), .A3(A[3]), .A4(n108), .Y(n76) );
  AO22X1_RVT U178 ( .A1(A_fpu[4]), .A2(n117), .A3(A[4]), .A4(n108), .Y(n77) );
  AO22X1_RVT U179 ( .A1(A_fpu[5]), .A2(n117), .A3(A[5]), .A4(n108), .Y(n78) );
  AO22X1_RVT U180 ( .A1(A_fpu[6]), .A2(n117), .A3(A[6]), .A4(n108), .Y(n79) );
  AO22X1_RVT U181 ( .A1(A_fpu[7]), .A2(n117), .A3(A[7]), .A4(n108), .Y(n80) );
  AO22X1_RVT U182 ( .A1(A_fpu[8]), .A2(n118), .A3(A[8]), .A4(n107), .Y(n81) );
  AO22X1_RVT U183 ( .A1(A_fpu[9]), .A2(n118), .A3(A[9]), .A4(n107), .Y(n82) );
  AO22X1_RVT U184 ( .A1(A_fpu[12]), .A2(n118), .A3(A[12]), .A4(n107), .Y(n85)
         );
  AO22X1_RVT U185 ( .A1(A_fpu[13]), .A2(n118), .A3(A[13]), .A4(n107), .Y(n86)
         );
  AO22X1_RVT U186 ( .A1(A_fpu[14]), .A2(n118), .A3(A[14]), .A4(n107), .Y(n87)
         );
  AO22X1_RVT U187 ( .A1(A_fpu[15]), .A2(n118), .A3(A[15]), .A4(n107), .Y(n88)
         );
  AO22X1_RVT U188 ( .A1(A_fpu[16]), .A2(n118), .A3(A[16]), .A4(n107), .Y(n89)
         );
  AO22X1_RVT U189 ( .A1(A_fpu[17]), .A2(n118), .A3(A[17]), .A4(n107), .Y(n90)
         );
  AO22X1_RVT U190 ( .A1(A_fpu[18]), .A2(n118), .A3(A[18]), .A4(n107), .Y(n91)
         );
  AO22X1_RVT U191 ( .A1(A_fpu[19]), .A2(n118), .A3(A[19]), .A4(n107), .Y(n92)
         );
  AO22X1_RVT U192 ( .A1(A_fpu[20]), .A2(n118), .A3(A[20]), .A4(n107), .Y(n93)
         );
  AO22X1_RVT U193 ( .A1(n111), .A2(Y[23]), .A3(Y_fpu[23]), .A4(n114), .Y(n14)
         );
  AO22X1_RVT U194 ( .A1(n111), .A2(Y[22]), .A3(Y_fpu[22]), .A4(n114), .Y(n15)
         );
  AO22X1_RVT U195 ( .A1(n111), .A2(Y[21]), .A3(Y_fpu[21]), .A4(n114), .Y(n16)
         );
  AO22X1_RVT U196 ( .A1(n111), .A2(Y[20]), .A3(Y_fpu[20]), .A4(n114), .Y(n17)
         );
  AO22X1_RVT U197 ( .A1(n111), .A2(Y[19]), .A3(Y_fpu[19]), .A4(n114), .Y(n18)
         );
  AO22X1_RVT U198 ( .A1(n111), .A2(Y[18]), .A3(Y_fpu[18]), .A4(n114), .Y(n19)
         );
  AO22X1_RVT U199 ( .A1(n111), .A2(Y[17]), .A3(Y_fpu[17]), .A4(n114), .Y(n20)
         );
  AO22X1_RVT U200 ( .A1(n111), .A2(Y[16]), .A3(Y_fpu[16]), .A4(n114), .Y(n21)
         );
  AO22X1_RVT U201 ( .A1(n111), .A2(Y[15]), .A3(Y_fpu[15]), .A4(n114), .Y(n22)
         );
  AO22X1_RVT U202 ( .A1(n105), .A2(n119), .A3(A[22]), .A4(n106), .Y(n95) );
  AO22X1_RVT U203 ( .A1(round_mode), .A2(n111), .A3(round_fpu), .A4(n114), .Y(
        n38) );
  INVX1_RVT U204 ( .A(start), .Y(n113) );
  INVX1_RVT U205 ( .A(reset), .Y(n127) );
  INVX1_RVT U206 ( .A(start), .Y(n115) );
  INVX1_RVT U207 ( .A(start), .Y(n117) );
  INVX1_RVT U208 ( .A(start), .Y(n116) );
  INVX1_RVT U209 ( .A(start), .Y(n118) );
  INVX1_RVT U210 ( .A(start), .Y(n114) );
  INVX1_RVT U211 ( .A(start), .Y(n119) );
  AO22X1_RVT U227 ( .A1(B_fpu[23]), .A2(n116), .A3(B[23]), .A4(n109), .Y(n64)
         );
  AO22X1_RVT U228 ( .A1(A_fpu[10]), .A2(n118), .A3(A[10]), .A4(n107), .Y(n83)
         );
  AO22X1_RVT U229 ( .A1(A_fpu[21]), .A2(n118), .A3(A[21]), .A4(n106), .Y(n94)
         );
endmodule
