`timescale 1ns/1ns
module tb_FPU;
reg Clock, Reset;
reg [31:0] A, B;
reg [1:0] Sel;
reg round;
reg start;
wire [31:0] Y;
wire Overflow, Error;

FPU FPU(Clock,Reset,A,B,Sel,round, start, Error,Overflow,Y);

initial
	$monitor($time, "A = %b, B = %b, Sel = %b, Y = %b, Overflow = %b, Error = %b", A, B, Sel, Y, Overflow, Error);

initial
begin
	Clock = 1'b0;
	forever #2 Clock = ~Clock;
end
	
initial begin 
	Reset=1;
	#3
	Reset=0;
	#2	
	Reset=1;
	A=32'b0_00010010_01101010100101000000000;
	B=32'b0_00001110_01110001001001000000000;
	Sel = 2'b00;
	start =1;
	round =0;
	#2
	start=0;
	#30

	A=32'b0_00010010_01101010100101000000000;
	B=32'b0_00001110_01110001001001000000000;
	Sel = 2'b00;
	start =1;
	round =1;
	#2
	start=0;
	#30

	A=32'b0_00010010_01101010100101000000000;
	B=32'b1_00001110_01110001001001000000000;
	Sel = 2'b00;
	start =1;
	round =0;
	#2
	start=0;
	#30

	A=32'b0_11111111_00000000000000000000000;
	B=32'b0_00001110_01110001001001000000000;
	Sel = 2'b00;
	start =1;
	round =0;
	#2
	start=0;
	#30

	A=32'b0_11111111_00000000000000000000000;
	B=32'b1_11111111_00000000000000000000000;
	Sel = 2'b00;
	start =1;
	round =0;
	#2
	start=0;
	#30

	A=32'b0_11111110_11100000000000000000000;
	B=32'b0_11111110_11100000000000000000000;
	Sel = 2'b00;
	start =1;
	round =0;
	#2
	start=0;
	#30

	A=32'b0_00000001_00001110000000000000000;
	B=32'b1_00000001_00000010110000000000000;
	Sel = 2'b00;
	start =1;
	round =0;
	#2
	start=0;
	#30

	A=32'b0_00010010_01101010100101000000000;
	B=32'b1_00001110_01110001001001000000000;
	Sel = 2'b01;
	start =1;
	round =0;
	#2
	start=0;
	#30

	A=32'b0_01010010_01100000000000000000000;
	B=32'b0_01001110_01110000000000000000000;
	Sel = 2'b10;
	start =1;
	round =0;
	#2
	start=0;
	#30

	A=32'b0_00010010_01100000000000000000000;
	B=32'b0_00001110_01110000000000000000000;
	Sel = 2'b10;
	start =1;
	round =0;
	#2
	start=0;
	#30

	A=32'b0_00010010_01100000000000000000000;
	B=32'b0_00000000_00000000000000000000000;
	Sel = 2'b10;
	start =1;
	round =0;
	#2
	start=0;
	#30

	A=32'b0_11111111_00000000000000000000000;
	B=32'b0_00001110_01110000000000000000000;
	Sel = 2'b10;
	start =1;
	round =0;
	#2
	start=0;
	#30

	A=32'b0_11111111_00000000000000000000000;
	B=32'b0_00000000_00000000000000000000000;
	Sel = 2'b10;
	start =1;
	round =0;
	#2
	start=0;
	#30

	A=32'b0_11111110_00000000000000000000000;
	B=32'b0_10000000_00000000000000000000000;
	Sel = 2'b10;
	start =1;
	round =0;
	#2
	start=0;
	#30

	A=32'b0_00001100_01000000000000000000000;
	B=32'b0_10000110_01000000000000000000000;
	Sel = 2'b11;
	start =1;
	round =0;
	#2
	start=0;
	#30

	A=32'b0_00001100_01000000000000000000000;
	B=32'b0_00000000_00000000000000000000000;
	Sel = 2'b11;
	start =1;
	round =0;
	#2
	start=0;
	#30

	A=32'b0_11111111_00000000000000000000000;
	B=32'b0_00000000_00000000000000000000000;
	Sel = 2'b11;
	start =1;
	round =0;
	#2
	start=0;
	#30

	A=32'b0_11111111_00000000000000000000000;
	B=32'b0_11111111_00000000000000000000000;
	Sel = 2'b11;
	start =1;
	round =0;
	#2
	start=0;
	#30

	A=32'b0_00000000_00000000000000000000000;
	B=32'b0_00000000_00000000000000000000000;
	Sel = 2'b11;
	start =1;
	round =0;
	#2
	start=0;
	#30

	A=32'b0_00001100_01000000000000000000000;
	B=32'b0_11111111_00000000000000000000000;
	Sel = 2'b11;
	start =1;
	round =0;
	#2
	start=0;
	#30

	A=32'b0_00000001_01000000000000000000000;
	B=32'b0_10000000_00000000000000000000000;
	Sel = 2'b11;
	start =1;
	round =0;
	#2
	start=0;
	#30
	$stop;
end

endmodule